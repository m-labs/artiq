/* Machine-generated using Migen */
module top(
	input serial_rx,
	output reg serial_tx,
	input clk125_gtp_p,
	input clk125_gtp_n,
	output [14:0] ddram_a,
	output [2:0] ddram_ba,
	output ddram_ras_n,
	output ddram_cas_n,
	output ddram_we_n,
	output [1:0] ddram_dm,
	inout [15:0] ddram_dq,
	output [1:0] ddram_dqs_p,
	output [1:0] ddram_dqs_n,
	output ddram_clk_p,
	output ddram_clk_n,
	output ddram_cke,
	output ddram_odt,
	output ddram_reset_n,
	output reg spiflash2x_cs_n,
	inout [1:0] spiflash2x_dq,
	input spiflash2x_wp,
	input spiflash2x_hold,
	output sfp_txp,
	output sfp_txn,
	input sfp_rxp,
	input sfp_rxn,
	output error_led,
	input cdr_clk_clean_p,
	input cdr_clk_clean_n,
	input sma_clkin_p,
	input sma_clkin_n,
	output cdr_clk_p,
	output cdr_clk_n,
	inout i2c_scl,
	inout i2c_sda,
	inout dio0_p,
	inout dio0_n,
	inout dio0_p_1,
	inout dio0_n_1,
	inout dio0_p_2,
	inout dio0_n_2,
	inout dio0_p_3,
	inout dio0_n_3,
	inout dio0_p_4,
	inout dio0_n_4,
	inout dio0_p_5,
	inout dio0_n_5,
	inout dio0_p_6,
	inout dio0_n_6,
	inout dio0_p_7,
	inout dio0_n_7,
	inout dio1_p,
	inout dio1_n,
	inout dio1_p_1,
	inout dio1_n_1,
	inout dio1_p_2,
	inout dio1_n_2,
	inout dio1_p_3,
	inout dio1_n_3,
	inout dio1_p_4,
	inout dio1_n_4,
	inout dio1_p_5,
	inout dio1_n_5,
	inout dio1_p_6,
	inout dio1_n_6,
	inout dio1_p_7,
	inout dio1_n_7,
	output urukul2_spi_p_clk,
	inout urukul2_spi_p_mosi,
	inout urukul2_spi_p_miso,
	output [2:0] urukul2_spi_p_cs_n,
	output urukul2_spi_n_clk,
	inout urukul2_spi_n_mosi,
	inout urukul2_spi_n_miso,
	output [2:0] urukul2_spi_n_cs_n,
	input urukul2_dds_reset_sync_in_p,
	input urukul2_dds_reset_sync_in_n,
	inout urukul2_io_update_p,
	inout urukul2_io_update_n,
	inout urukul2_sw0_p,
	inout urukul2_sw0_n,
	inout urukul2_sw1_p,
	inout urukul2_sw1_n,
	inout urukul2_sw2_p,
	inout urukul2_sw2_n,
	inout urukul2_sw3_p,
	inout urukul2_sw3_n,
	output urukul4_spi_p_clk,
	inout urukul4_spi_p_mosi,
	inout urukul4_spi_p_miso,
	output [2:0] urukul4_spi_p_cs_n,
	output urukul4_spi_n_clk,
	inout urukul4_spi_n_mosi,
	inout urukul4_spi_n_miso,
	output [2:0] urukul4_spi_n_cs_n,
	output urukul4_dds_reset_sync_in_p,
	output urukul4_dds_reset_sync_in_n,
	inout urukul4_io_update_p,
	inout urukul4_io_update_n,
	inout urukul4_sw0_p,
	inout urukul4_sw0_n,
	inout urukul4_sw1_p,
	inout urukul4_sw1_n,
	inout urukul4_sw2_p,
	inout urukul4_sw2_n,
	inout urukul4_sw3_p,
	inout urukul4_sw3_n,
	output sampler6_adc_spi_p_clk,
	inout sampler6_adc_spi_p_miso,
	output sampler6_adc_spi_n_clk,
	inout sampler6_adc_spi_n_miso,
	output sampler6_pgia_spi_p_clk,
	inout sampler6_pgia_spi_p_mosi,
	inout sampler6_pgia_spi_p_miso,
	output sampler6_pgia_spi_p_cs_n,
	output sampler6_pgia_spi_n_clk,
	inout sampler6_pgia_spi_n_mosi,
	inout sampler6_pgia_spi_n_miso,
	output sampler6_pgia_spi_n_cs_n,
	inout sampler6_cnv_p,
	inout sampler6_cnv_n,
	output sampler6_sdr_p,
	output sampler6_sdr_n,
	output zotino8_spi_p_clk,
	inout zotino8_spi_p_mosi,
	inout zotino8_spi_p_miso,
	output [1:0] zotino8_spi_p_cs_n,
	output zotino8_spi_n_clk,
	inout zotino8_spi_n_mosi,
	inout zotino8_spi_n_miso,
	output [1:0] zotino8_spi_n_cs_n,
	inout zotino8_ldac_n_p,
	inout zotino8_ldac_n_n,
	inout zotino8_clr_n_p,
	inout zotino8_clr_n_n,
	output user_led,
	output user_led_1,
	output user_led_2
);

wire [28:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_adr;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_w;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_bte;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_err;
wire [28:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_adr;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_w;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_dbus_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_dbus_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_dbus_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_dbus_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_bte;
wire main_genericstandalone_genericstandalone_genericstandalone_dbus_err;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_interrupt;
wire [28:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_adr;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_w;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_sram_bus_err = 1'd0;
wire [9:0] main_genericstandalone_genericstandalone_genericstandalone_sram_adr;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_sram_dat_r;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_sram_we;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w;
reg [13:0] main_genericstandalone_genericstandalone_genericstandalone_interface_adr = 14'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_interface_we = 1'd0;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w = 8'd0;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_interface_dat_r;
wire [28:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_adr;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_w;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_r = 64'd0;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_err = 1'd0;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_trigger = 2'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full = 32'd3958241;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_last;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_payload_data;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx = 32'd0;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg = 8'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount = 4'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_ack;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_last = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_eop = 1'd0;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_payload_data = 8'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx = 32'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_r = 1'd0;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg = 8'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount = 4'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_re;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_w;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_txfull_status;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rxempty_status;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_irq;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_status;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_clear;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_old_trigger = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_status;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_rx_old_trigger = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_status_re;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_status_r;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_status_w;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_pending_re;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_pending_r;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full = 2'd0;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_ack;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_eop = 1'd0;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_ack;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_last = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_re;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_readable;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_din;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_dout;
reg [4:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level = 5'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce = 4'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume = 4'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_r;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_we;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_w;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_adr;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_eop;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_last;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_re;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_readable;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_din;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_dout;
reg [4:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level = 5'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce = 4'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume = 4'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_r;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_we;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_w;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_adr;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_eop;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full = 64'd0;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_load_re = 1'd0;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full = 64'd0;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_re = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_en_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_re;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_r;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_w = 1'd0;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status = 64'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_irq;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_status;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_clear;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_old_trigger = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_re;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_r;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_w;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_re;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_r;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_w;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_re = 1'd0;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_value = 64'd0;
wire [28:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_w;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_err = 1'd0;
wire sys_clk;
wire sys_rst;
wire sys4x_clk;
wire sys4x_dqs_clk;
wire clk200_clk;
wire clk200_rst;
wire bootstrap_clk;
wire main_genericstandalone_genericstandalone_crg_status;
wire main_genericstandalone_genericstandalone_crg_clk125_buf;
wire main_genericstandalone_genericstandalone_crg_clk125_div2_raw;
wire main_genericstandalone_genericstandalone_crg_clk125_div2;
(* dont_touch = "true" *) wire main_genericstandalone_genericstandalone_crg_i_clk_sw;
(* dont_touch = "true" *) reg main_genericstandalone_genericstandalone_crg_o_clk_sw = 1'd0;
(* dont_touch = "true" *) reg main_genericstandalone_genericstandalone_crg_o_reset = 1'd0;
(* dont_touch = "true" *) wire main_genericstandalone_genericstandalone_crg_i_switch;
reg main_genericstandalone_genericstandalone_crg_o_switch = 1'd0;
reg main_genericstandalone_genericstandalone_crg_reset;
reg [15:0] main_genericstandalone_genericstandalone_crg_delay_counter = 16'd65535;
wire main_genericstandalone_genericstandalone_crg_pll_clk200;
wire main_genericstandalone_genericstandalone_crg_pll_clk_bootstrap;
wire main_genericstandalone_genericstandalone_crg_pll_fb;
wire main_genericstandalone_genericstandalone_crg_pll_locked;
reg [3:0] main_genericstandalone_genericstandalone_crg_reset_counter = 4'd15;
reg main_genericstandalone_genericstandalone_crg_ic_reset = 1'd1;
reg [1:0] main_genericstandalone_genericstandalone_ddrphy_storage_full = 2'd0;
wire [1:0] main_genericstandalone_genericstandalone_ddrphy_storage;
reg main_genericstandalone_genericstandalone_ddrphy_re = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_r;
reg main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_w = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_r;
reg main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_w = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_r;
reg main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_w = 1'd0;
wire [14:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address;
wire [2:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cas_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cs_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_ras_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_we_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cke;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_odt;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata;
reg main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_valid = 1'd0;
wire [14:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address;
wire [2:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cas_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cs_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_ras_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_we_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cke;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_odt;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata;
reg main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_valid = 1'd0;
wire [14:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address;
wire [2:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cas_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cs_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_ras_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_we_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cke;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_odt;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata;
reg main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_valid = 1'd0;
wire [14:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address;
wire [2:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cas_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cs_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_ras_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_we_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cke;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_odt;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata;
reg main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_valid = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_sd_clk_se;
reg main_genericstandalone_genericstandalone_ddrphy_oe_dqs = 1'd0;
reg [7:0] main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern = 8'd85;
wire main_genericstandalone_genericstandalone_ddrphy_dqs0;
wire main_genericstandalone_genericstandalone_ddrphy_dqs_t0;
wire main_genericstandalone_genericstandalone_ddrphy_dqs1;
wire main_genericstandalone_genericstandalone_ddrphy_dqs_t1;
reg main_genericstandalone_genericstandalone_ddrphy_oe_dq = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o1;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay1;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed1;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t1;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o2;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay2;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed2;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t2;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o3;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay3;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed3;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t3;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o4;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay4;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed4;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t4;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o5;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay5;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed5;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t5;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o6;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay6;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed6;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t6;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o7;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay7;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed7;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t7;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o8;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay8;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed8;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t8;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o9;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay9;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed9;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t9;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o10;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay10;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed10;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t10;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o11;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay11;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed11;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t11;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o12;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay12;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed12;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t12;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o13;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay13;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed13;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t13;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o14;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay14;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed14;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t14;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o15;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay15;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed15;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t15;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en0 = 1'd0;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en1 = 1'd0;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en2 = 1'd0;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en3 = 1'd0;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4 = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_oe;
reg [3:0] main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en = 4'd0;
wire [28:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_adr;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_w;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_bte;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_err;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_bank;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cs_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_ras_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_bank;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cs_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_ras_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_bank;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cs_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_ras_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_bank;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cs_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_ras_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_address;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_address;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_address;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_address;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_valid;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_storage_full = 4'd0;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_re = 1'd0;
reg [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full = 6'd0;
wire [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_r;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_w = 1'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full = 15'd0;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_re = 1'd0;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full = 3'd0;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full = 32'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status = 32'd0;
reg [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full = 6'd0;
wire [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_r;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_w = 1'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full = 15'd0;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_re = 1'd0;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full = 3'd0;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full = 32'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status = 32'd0;
reg [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full = 6'd0;
wire [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_r;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_w = 1'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full = 15'd0;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_re = 1'd0;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full = 3'd0;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full = 32'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status = 32'd0;
reg [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full = 6'd0;
wire [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_r;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_w = 1'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full = 15'd0;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_re = 1'd0;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full = 3'd0;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full = 32'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status = 32'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata = 32'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_en = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_mask = 4'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata_en = 1'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata = 32'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_en = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_mask = 4'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata = 32'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_mask = 4'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata_en = 1'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cas_n = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_ras_n = 1'd1;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_we_n = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata = 32'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_en = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_mask = 4'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata_en = 1'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata_valid;
wire [28:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_w;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r;
wire [15:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_err = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_idle;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_hit;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset0;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset2;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset3;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset4;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset5;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset6;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset7;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_wait;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_done;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_count = 3'd4;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_pending_refresh = 1'd0;
reg [9:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refi_cycles = 10'd977;
reg [9:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col = 10'd0;
wire [9:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col_inc_next;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_swap_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_adr_inc;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_burst;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_rdvalid_r = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read_ended;
reg [127:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_dat_w0 = 128'd0;
reg [15:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_sel0 = 16'd0;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_dat_w1;
wire [15:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_sel1;
wire [28:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_adr;
reg [127:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_r;
wire [15:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_sel;
reg main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc;
reg main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack;
reg main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cti;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_bte = 2'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_err;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_cache = 2'd0;
wire [10:0] main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_adr;
wire [511:0] main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_we;
reg [511:0] main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_w;
reg main_genericstandalone_genericstandalone_genericstandalone_cache_write_from_slave;
reg main_genericstandalone_genericstandalone_genericstandalone_cache_adr_inc;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_cache_next_adr_offset;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_cache_adr_offset_r = 3'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_cache_last;
wire main_genericstandalone_genericstandalone_genericstandalone_cache_newline;
wire [10:0] main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_adr;
wire [16:0] main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_dat_r;
reg main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_we;
wire [16:0] main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_dat_w;
wire [15:0] main_genericstandalone_genericstandalone_genericstandalone_cache_tag_do_tag;
wire main_genericstandalone_genericstandalone_genericstandalone_cache_tag_do_dirty;
wire [15:0] main_genericstandalone_genericstandalone_genericstandalone_cache_tag_di_tag;
reg main_genericstandalone_genericstandalone_genericstandalone_cache_tag_di_dirty;
reg main_genericstandalone_genericstandalone_genericstandalone_cache_word_clr;
reg main_genericstandalone_genericstandalone_genericstandalone_cache_word_inc;
wire [7:0] main_genericstandalone_genericstandalone_virtual_leds_status;
reg main_genericstandalone_genericstandalone_clk;
wire [28:0] main_genericstandalone_genericstandalone_spiflash_bus_adr;
wire [63:0] main_genericstandalone_genericstandalone_spiflash_bus_dat_w;
wire [63:0] main_genericstandalone_genericstandalone_spiflash_bus_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_spiflash_bus_sel;
wire main_genericstandalone_genericstandalone_spiflash_bus_cyc;
wire main_genericstandalone_genericstandalone_spiflash_bus_stb;
reg main_genericstandalone_genericstandalone_spiflash_bus_ack = 1'd0;
wire main_genericstandalone_genericstandalone_spiflash_bus_we;
wire [2:0] main_genericstandalone_genericstandalone_spiflash_bus_cti;
wire [1:0] main_genericstandalone_genericstandalone_spiflash_bus_bte;
reg main_genericstandalone_genericstandalone_spiflash_bus_err = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full = 4'd0;
wire [3:0] main_genericstandalone_genericstandalone_spiflash_bitbang_storage;
reg main_genericstandalone_genericstandalone_spiflash_bitbang_re = 1'd0;
reg main_genericstandalone_genericstandalone_spiflash_status;
reg main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full = 1'd0;
wire main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage;
reg main_genericstandalone_genericstandalone_spiflash_bitbang_en_re = 1'd0;
reg main_genericstandalone_genericstandalone_spiflash_cs_n = 1'd1;
reg main_genericstandalone_genericstandalone_spiflash_clk = 1'd0;
reg main_genericstandalone_genericstandalone_spiflash_dq_oe = 1'd0;
reg [1:0] main_genericstandalone_genericstandalone_spiflash_o;
reg main_genericstandalone_genericstandalone_spiflash_oe;
wire [1:0] main_genericstandalone_genericstandalone_spiflash_i0;
reg [63:0] main_genericstandalone_genericstandalone_spiflash_sr = 64'd0;
reg main_genericstandalone_genericstandalone_spiflash_i1 = 1'd0;
reg [1:0] main_genericstandalone_genericstandalone_spiflash_dqi = 2'd0;
reg [6:0] main_genericstandalone_genericstandalone_spiflash_trigger = 7'd0;
wire main_genericstandalone_genericstandalone_icap_iprog_re;
wire main_genericstandalone_genericstandalone_icap_iprog_r;
reg main_genericstandalone_genericstandalone_icap_iprog_w = 1'd0;
reg main_genericstandalone_genericstandalone_icap_icap_csib;
reg [31:0] main_genericstandalone_genericstandalone_icap_icap_i;
reg main_genericstandalone_genericstandalone_icap_icap_rdwrb;
wire icap_clk;
reg main_genericstandalone_genericstandalone_icap_counter0 = 1'd0;
wire main_genericstandalone_genericstandalone_icap_counter_rst;
wire main_genericstandalone_genericstandalone_icap_i;
wire main_genericstandalone_genericstandalone_icap_o;
reg main_genericstandalone_genericstandalone_icap_toggle_i = 1'd0;
wire main_genericstandalone_genericstandalone_icap_toggle_o;
reg main_genericstandalone_genericstandalone_icap_toggle_o_r = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_icap_counter1 = 4'd0;
wire main_genericstandalone_genericstandalone_qpll_reset;
wire main_genericstandalone_genericstandalone_qpll_lock;
wire main_genericstandalone_genericstandalone_qpll_clk;
wire main_genericstandalone_genericstandalone_qpll_refclk;
reg main_genericstandalone_pcs_transmitpath_config_stb;
wire [15:0] main_genericstandalone_pcs_transmitpath_config_reg;
wire main_genericstandalone_pcs_transmitpath_tx_stb;
reg main_genericstandalone_pcs_transmitpath_tx_ack;
wire [7:0] main_genericstandalone_pcs_transmitpath_tx_data;
reg [7:0] main_genericstandalone_pcs_transmitpath_encoder0;
reg main_genericstandalone_pcs_transmitpath_encoder1;
reg [9:0] main_genericstandalone_pcs_transmitpath_encoder2 = 10'd0;
reg main_genericstandalone_pcs_transmitpath_encoder3 = 1'd0;
wire [7:0] main_genericstandalone_pcs_transmitpath_encoder_d;
wire main_genericstandalone_pcs_transmitpath_encoder_k;
reg main_genericstandalone_pcs_transmitpath_encoder_disp_in = 1'd0;
reg [9:0] main_genericstandalone_pcs_transmitpath_encoder_output;
reg main_genericstandalone_pcs_transmitpath_encoder_disp_out;
reg [5:0] main_genericstandalone_pcs_transmitpath_encoder_code6b = 6'd0;
reg main_genericstandalone_pcs_transmitpath_encoder_code6b_unbalanced = 1'd0;
reg main_genericstandalone_pcs_transmitpath_encoder_code6b_flip = 1'd0;
reg [3:0] main_genericstandalone_pcs_transmitpath_encoder_code4b = 4'd0;
reg main_genericstandalone_pcs_transmitpath_encoder_code4b_unbalanced = 1'd0;
reg main_genericstandalone_pcs_transmitpath_encoder_code4b_flip = 1'd0;
reg main_genericstandalone_pcs_transmitpath_encoder_alt7_rd0 = 1'd0;
reg main_genericstandalone_pcs_transmitpath_encoder_alt7_rd1 = 1'd0;
reg [5:0] main_genericstandalone_pcs_transmitpath_encoder_output_6b;
wire main_genericstandalone_pcs_transmitpath_encoder_disp_inter;
reg [3:0] main_genericstandalone_pcs_transmitpath_encoder_output_4b;
wire [9:0] main_genericstandalone_pcs_transmitpath_encoder_output_msb_first;
wire [1:0] main_genericstandalone_pcs_transmitpath_sgmii_speed;
reg main_genericstandalone_pcs_transmitpath_parity = 1'd0;
reg main_genericstandalone_pcs_transmitpath_c_type = 1'd0;
reg [15:0] main_genericstandalone_pcs_transmitpath_config_reg_buffer = 16'd0;
reg main_genericstandalone_pcs_transmitpath_load_config_reg_buffer;
reg [9:0] main_genericstandalone_pcs_transmitpath_timer = 10'd0;
reg main_genericstandalone_pcs_transmitpath_timer_en;
reg main_genericstandalone_pcs_receivepath_rx_en;
wire [7:0] main_genericstandalone_pcs_receivepath_rx_data;
reg main_genericstandalone_pcs_receivepath_seen_valid_ci;
reg main_genericstandalone_pcs_receivepath_seen_config_reg = 1'd0;
reg [15:0] main_genericstandalone_pcs_receivepath_config_reg = 16'd0;
wire [9:0] main_genericstandalone_pcs_receivepath_input;
wire [7:0] main_genericstandalone_pcs_receivepath_d;
reg main_genericstandalone_pcs_receivepath_k = 1'd0;
reg [9:0] main_genericstandalone_pcs_receivepath_input_msb_first;
reg [4:0] main_genericstandalone_pcs_receivepath_code5b = 5'd0;
reg [2:0] main_genericstandalone_pcs_receivepath_code3b = 3'd0;
wire [1:0] main_genericstandalone_pcs_receivepath_sgmii_speed;
wire main_genericstandalone_pcs_receivepath_sample_en;
reg [7:0] main_genericstandalone_pcs_receivepath_config_reg_lsb = 8'd0;
reg main_genericstandalone_pcs_receivepath_load_config_reg_lsb;
reg main_genericstandalone_pcs_receivepath_load_config_reg_msb;
reg main_genericstandalone_pcs_receivepath_first_preamble_byte;
reg [9:0] main_genericstandalone_pcs_receivepath_timer = 10'd0;
reg main_genericstandalone_pcs_receivepath_timer_en;
wire main_genericstandalone_pcs_sink_stb;
wire main_genericstandalone_pcs_sink_ack;
wire main_genericstandalone_pcs_sink_last;
wire main_genericstandalone_pcs_sink_eop;
wire [7:0] main_genericstandalone_pcs_sink_payload_data;
wire main_genericstandalone_pcs_sink_payload_last_be;
wire main_genericstandalone_pcs_sink_payload_error;
reg main_genericstandalone_pcs_source_stb = 1'd0;
wire main_genericstandalone_pcs_source_ack;
reg main_genericstandalone_pcs_source_last = 1'd0;
wire main_genericstandalone_pcs_source_eop;
reg [7:0] main_genericstandalone_pcs_source_payload_data = 8'd0;
reg main_genericstandalone_pcs_source_payload_last_be = 1'd0;
reg main_genericstandalone_pcs_source_payload_error = 1'd0;
reg main_genericstandalone_pcs_link_up;
reg main_genericstandalone_pcs_restart;
reg [15:0] main_genericstandalone_pcs_lp_abi_i = 16'd0;
reg [15:0] main_genericstandalone_pcs_lp_abi_o = 16'd0;
reg main_genericstandalone_pcs_lp_abi_starter = 1'd1;
wire main_genericstandalone_pcs_lp_abi_ping_i;
wire main_genericstandalone_pcs_lp_abi_ping_o0;
reg main_genericstandalone_pcs_lp_abi_ping_toggle_i = 1'd0;
wire main_genericstandalone_pcs_lp_abi_ping_toggle_o;
reg main_genericstandalone_pcs_lp_abi_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_pcs_lp_abi_ping_o1 = 1'd0;
wire main_genericstandalone_pcs_lp_abi_pong_i;
wire main_genericstandalone_pcs_lp_abi_pong_o;
reg main_genericstandalone_pcs_lp_abi_pong_toggle_i = 1'd0;
wire main_genericstandalone_pcs_lp_abi_pong_toggle_o;
reg main_genericstandalone_pcs_lp_abi_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_pcs_lp_abi_wait;
wire main_genericstandalone_pcs_lp_abi_done;
reg [7:0] main_genericstandalone_pcs_lp_abi_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_pcs_lp_abi_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_pcs_lp_abi_obuffer;
reg main_genericstandalone_pcs_rx_en_d = 1'd0;
wire main_genericstandalone_pcs_seen_valid_ci_i;
wire main_genericstandalone_pcs_seen_valid_ci_o;
reg main_genericstandalone_pcs_seen_valid_ci_toggle_i = 1'd0;
wire main_genericstandalone_pcs_seen_valid_ci_toggle_o;
reg main_genericstandalone_pcs_seen_valid_ci_toggle_o_r = 1'd0;
reg [19:0] main_genericstandalone_pcs_checker_counter = 20'd0;
reg main_genericstandalone_pcs_checker_tick = 1'd0;
reg main_genericstandalone_pcs_checker_ok = 1'd0;
reg main_genericstandalone_pcs_tx_config_empty;
wire main_genericstandalone_pcs_is_sgmii;
wire main_genericstandalone_pcs_linkdown;
reg main_genericstandalone_pcs_autoneg_ack;
reg main_genericstandalone_pcs_rx_config_reg_abi_i = 1'd0;
wire main_genericstandalone_pcs_rx_config_reg_abi_o;
reg main_genericstandalone_pcs_rx_config_reg_abi_toggle_i = 1'd0;
wire main_genericstandalone_pcs_rx_config_reg_abi_toggle_o;
reg main_genericstandalone_pcs_rx_config_reg_abi_toggle_o_r = 1'd0;
reg main_genericstandalone_pcs_rx_config_reg_ack_i = 1'd0;
wire main_genericstandalone_pcs_rx_config_reg_ack_o;
reg main_genericstandalone_pcs_rx_config_reg_ack_toggle_i = 1'd0;
wire main_genericstandalone_pcs_rx_config_reg_ack_toggle_o;
reg main_genericstandalone_pcs_rx_config_reg_ack_toggle_o_r = 1'd0;
reg main_genericstandalone_pcs_waittimer0_wait;
wire main_genericstandalone_pcs_waittimer0_done;
reg [20:0] main_genericstandalone_pcs_waittimer0_count = 21'd1250000;
reg main_genericstandalone_pcs_waittimer1_wait;
wire main_genericstandalone_pcs_waittimer1_done;
reg [17:0] main_genericstandalone_pcs_waittimer1_count = 18'd200000;
reg [2:0] main_genericstandalone_pcs_c_counter = 3'd0;
reg [15:0] main_genericstandalone_pcs_prev_config_reg = 16'd0;
wire eth_tx_clk;
wire eth_tx_rst;
wire eth_rx_clk;
wire eth_rx_rst;
wire eth_tx_half_clk;
wire eth_rx_half_clk;
wire main_genericstandalone_txoutclk;
wire main_genericstandalone_rxoutclk;
wire main_genericstandalone_tx_reset;
wire main_genericstandalone_tx_mmcm_locked;
wire [19:0] main_genericstandalone_tx_data0;
wire main_genericstandalone_tx_reset_done;
wire main_genericstandalone_rx_reset;
wire main_genericstandalone_rx_mmcm_locked;
wire [19:0] main_genericstandalone_rx_data0;
wire main_genericstandalone_rx_reset_done;
wire main_genericstandalone_rx_pma_reset_done;
wire [8:0] main_genericstandalone_drpaddr;
wire main_genericstandalone_drpen;
wire [15:0] main_genericstandalone_drpdi;
wire main_genericstandalone_drprdy;
wire [15:0] main_genericstandalone_drpdo;
wire main_genericstandalone_drpwe;
wire main_genericstandalone_txoutclk_rebuffer;
wire main_genericstandalone_rxoutclk_rebuffer;
wire main_genericstandalone_tx_mmcm_fb;
(* dont_touch = "true" *) reg main_genericstandalone_tx_mmcm_reset = 1'd1;
wire main_genericstandalone_clk_tx_unbuf;
wire main_genericstandalone_clk_tx_half_unbuf;
wire main_genericstandalone_rx_mmcm_fb;
(* dont_touch = "true" *) reg main_genericstandalone_rx_mmcm_reset = 1'd1;
wire main_genericstandalone_clk_rx_unbuf;
wire main_genericstandalone_clk_rx_half_unbuf;
(* dont_touch = "true" *) reg main_genericstandalone_tx_init_qpll_reset0 = 1'd0;
wire main_genericstandalone_tx_init_qpll_lock0;
(* dont_touch = "true" *) reg main_genericstandalone_tx_init_tx_reset0 = 1'd0;
reg main_genericstandalone_tx_init_done;
reg main_genericstandalone_tx_init_qpll_reset1;
reg main_genericstandalone_tx_init_tx_reset1;
wire main_genericstandalone_tx_init_qpll_lock1;
reg [5:0] main_genericstandalone_tx_init_timer = 6'd0;
reg main_genericstandalone_tx_init_tick = 1'd0;
(* dont_touch = "true" *) reg main_genericstandalone_rx_init_rx_reset0 = 1'd0;
wire main_genericstandalone_rx_init_rx_pma_reset_done0;
wire [8:0] main_genericstandalone_rx_init_drpaddr;
reg main_genericstandalone_rx_init_drpen;
reg [15:0] main_genericstandalone_rx_init_drpdi;
wire main_genericstandalone_rx_init_drprdy;
wire [15:0] main_genericstandalone_rx_init_drpdo;
reg main_genericstandalone_rx_init_drpwe;
wire main_genericstandalone_rx_init_enable;
wire main_genericstandalone_rx_init_restart;
reg main_genericstandalone_rx_init_done;
reg main_genericstandalone_rx_init_rx_reset1;
wire main_genericstandalone_rx_init_rx_pma_reset_done1;
reg [15:0] main_genericstandalone_rx_init_drpvalue = 16'd0;
reg main_genericstandalone_rx_init_drpmask;
reg main_genericstandalone_rx_init_rx_pma_reset_done_r = 1'd0;
wire main_genericstandalone_i;
wire main_genericstandalone_o;
reg main_genericstandalone_toggle_i = 1'd0;
wire main_genericstandalone_toggle_o;
reg main_genericstandalone_toggle_o_r = 1'd0;
reg [12:0] main_genericstandalone_cdr_lock_counter = 13'd0;
reg main_genericstandalone_cdr_locked = 1'd0;
wire [9:0] main_genericstandalone_tx_data1;
reg [19:0] main_genericstandalone_tx_data_half = 20'd0;
wire [19:0] main_genericstandalone_rx_data_half;
reg [9:0] main_genericstandalone_rx_data1 = 10'd0;
reg [19:0] main_genericstandalone_buf = 20'd0;
reg main_genericstandalone_phase_half = 1'd0;
reg main_genericstandalone_phase_half_rereg = 1'd0;
wire main_genericstandalone_virtual_led;
wire main_genericstandalone_tx_gap_inserter_sink_stb;
reg main_genericstandalone_tx_gap_inserter_sink_ack;
wire main_genericstandalone_tx_gap_inserter_sink_last;
wire main_genericstandalone_tx_gap_inserter_sink_eop;
wire [7:0] main_genericstandalone_tx_gap_inserter_sink_payload_data;
wire main_genericstandalone_tx_gap_inserter_sink_payload_last_be;
wire main_genericstandalone_tx_gap_inserter_sink_payload_error;
reg main_genericstandalone_tx_gap_inserter_source_stb;
wire main_genericstandalone_tx_gap_inserter_source_ack;
reg main_genericstandalone_tx_gap_inserter_source_last;
reg main_genericstandalone_tx_gap_inserter_source_eop;
reg [7:0] main_genericstandalone_tx_gap_inserter_source_payload_data;
reg main_genericstandalone_tx_gap_inserter_source_payload_last_be;
reg main_genericstandalone_tx_gap_inserter_source_payload_error;
reg [3:0] main_genericstandalone_tx_gap_inserter_counter = 4'd0;
reg main_genericstandalone_tx_gap_inserter_counter_reset;
reg main_genericstandalone_tx_gap_inserter_counter_ce;
reg [31:0] main_genericstandalone_preamble_errors_status = 32'd0;
reg [31:0] main_genericstandalone_crc_errors_status = 32'd0;
wire main_genericstandalone_preamble_inserter_sink_stb;
reg main_genericstandalone_preamble_inserter_sink_ack;
wire main_genericstandalone_preamble_inserter_sink_last;
wire main_genericstandalone_preamble_inserter_sink_eop;
wire [7:0] main_genericstandalone_preamble_inserter_sink_payload_data;
wire main_genericstandalone_preamble_inserter_sink_payload_last_be;
wire main_genericstandalone_preamble_inserter_sink_payload_error;
reg main_genericstandalone_preamble_inserter_source_stb;
wire main_genericstandalone_preamble_inserter_source_ack;
reg main_genericstandalone_preamble_inserter_source_last;
reg main_genericstandalone_preamble_inserter_source_eop;
reg [7:0] main_genericstandalone_preamble_inserter_source_payload_data;
wire main_genericstandalone_preamble_inserter_source_payload_last_be;
reg main_genericstandalone_preamble_inserter_source_payload_error;
reg [63:0] main_genericstandalone_preamble_inserter_preamble = 64'd15372286728091293013;
reg [2:0] main_genericstandalone_preamble_inserter_cnt = 3'd0;
reg main_genericstandalone_preamble_inserter_clr_cnt;
reg main_genericstandalone_preamble_inserter_inc_cnt;
wire main_genericstandalone_preamble_checker_sink_stb;
reg main_genericstandalone_preamble_checker_sink_ack;
wire main_genericstandalone_preamble_checker_sink_last;
wire main_genericstandalone_preamble_checker_sink_eop;
wire [7:0] main_genericstandalone_preamble_checker_sink_payload_data;
wire main_genericstandalone_preamble_checker_sink_payload_last_be;
wire main_genericstandalone_preamble_checker_sink_payload_error;
reg main_genericstandalone_preamble_checker_source_stb;
wire main_genericstandalone_preamble_checker_source_ack;
reg main_genericstandalone_preamble_checker_source_last;
reg main_genericstandalone_preamble_checker_source_eop;
wire [7:0] main_genericstandalone_preamble_checker_source_payload_data;
wire main_genericstandalone_preamble_checker_source_payload_last_be;
reg main_genericstandalone_preamble_checker_source_payload_error;
reg main_genericstandalone_preamble_checker_error;
wire main_genericstandalone_crc32_inserter_sink_stb;
reg main_genericstandalone_crc32_inserter_sink_ack;
wire main_genericstandalone_crc32_inserter_sink_last;
wire main_genericstandalone_crc32_inserter_sink_eop;
wire [7:0] main_genericstandalone_crc32_inserter_sink_payload_data;
wire main_genericstandalone_crc32_inserter_sink_payload_last_be;
wire main_genericstandalone_crc32_inserter_sink_payload_error;
reg main_genericstandalone_crc32_inserter_source_stb;
wire main_genericstandalone_crc32_inserter_source_ack;
reg main_genericstandalone_crc32_inserter_source_last;
reg main_genericstandalone_crc32_inserter_source_eop;
reg [7:0] main_genericstandalone_crc32_inserter_source_payload_data;
reg main_genericstandalone_crc32_inserter_source_payload_last_be;
reg main_genericstandalone_crc32_inserter_source_payload_error;
reg [7:0] main_genericstandalone_crc32_inserter_data0;
wire [31:0] main_genericstandalone_crc32_inserter_value;
wire main_genericstandalone_crc32_inserter_error;
wire [7:0] main_genericstandalone_crc32_inserter_data1;
wire [31:0] main_genericstandalone_crc32_inserter_last;
reg [31:0] main_genericstandalone_crc32_inserter_next;
reg [31:0] main_genericstandalone_crc32_inserter_reg = 32'd4294967295;
reg main_genericstandalone_crc32_inserter_ce;
reg main_genericstandalone_crc32_inserter_reset;
reg [1:0] main_genericstandalone_crc32_inserter_cnt = 2'd3;
wire main_genericstandalone_crc32_inserter_cnt_done;
reg main_genericstandalone_crc32_inserter_is_ongoing0;
reg main_genericstandalone_crc32_inserter_is_ongoing1;
wire main_genericstandalone_crc32_checker_sink_sink_stb;
reg main_genericstandalone_crc32_checker_sink_sink_ack;
wire main_genericstandalone_crc32_checker_sink_sink_last;
wire main_genericstandalone_crc32_checker_sink_sink_eop;
wire [7:0] main_genericstandalone_crc32_checker_sink_sink_payload_data;
wire main_genericstandalone_crc32_checker_sink_sink_payload_last_be;
wire main_genericstandalone_crc32_checker_sink_sink_payload_error;
wire main_genericstandalone_crc32_checker_source_source_stb;
wire main_genericstandalone_crc32_checker_source_source_ack;
reg main_genericstandalone_crc32_checker_source_source_last = 1'd0;
wire main_genericstandalone_crc32_checker_source_source_eop;
wire [7:0] main_genericstandalone_crc32_checker_source_source_payload_data;
wire main_genericstandalone_crc32_checker_source_source_payload_last_be;
reg main_genericstandalone_crc32_checker_source_source_payload_error;
wire main_genericstandalone_crc32_checker_error;
wire [7:0] main_genericstandalone_crc32_checker_crc_data0;
wire [31:0] main_genericstandalone_crc32_checker_crc_value;
wire main_genericstandalone_crc32_checker_crc_error;
wire [7:0] main_genericstandalone_crc32_checker_crc_data1;
wire [31:0] main_genericstandalone_crc32_checker_crc_last;
reg [31:0] main_genericstandalone_crc32_checker_crc_next;
reg [31:0] main_genericstandalone_crc32_checker_crc_reg = 32'd4294967295;
reg main_genericstandalone_crc32_checker_crc_ce;
reg main_genericstandalone_crc32_checker_crc_reset;
reg main_genericstandalone_crc32_checker_syncfifo_sink_stb;
wire main_genericstandalone_crc32_checker_syncfifo_sink_ack;
wire main_genericstandalone_crc32_checker_syncfifo_sink_last;
wire main_genericstandalone_crc32_checker_syncfifo_sink_eop;
wire [7:0] main_genericstandalone_crc32_checker_syncfifo_sink_payload_data;
wire main_genericstandalone_crc32_checker_syncfifo_sink_payload_last_be;
wire main_genericstandalone_crc32_checker_syncfifo_sink_payload_error;
wire main_genericstandalone_crc32_checker_syncfifo_source_stb;
wire main_genericstandalone_crc32_checker_syncfifo_source_ack;
wire main_genericstandalone_crc32_checker_syncfifo_source_eop;
wire [7:0] main_genericstandalone_crc32_checker_syncfifo_source_payload_data;
wire main_genericstandalone_crc32_checker_syncfifo_source_payload_last_be;
wire main_genericstandalone_crc32_checker_syncfifo_source_payload_error;
wire main_genericstandalone_crc32_checker_syncfifo_syncfifo_we;
wire main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable;
wire main_genericstandalone_crc32_checker_syncfifo_syncfifo_re;
wire main_genericstandalone_crc32_checker_syncfifo_syncfifo_readable;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_syncfifo_din;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_syncfifo_dout;
reg [2:0] main_genericstandalone_crc32_checker_syncfifo_level = 3'd0;
reg main_genericstandalone_crc32_checker_syncfifo_replace = 1'd0;
reg [2:0] main_genericstandalone_crc32_checker_syncfifo_produce = 3'd0;
reg [2:0] main_genericstandalone_crc32_checker_syncfifo_consume = 3'd0;
reg [2:0] main_genericstandalone_crc32_checker_syncfifo_wrport_adr;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_wrport_dat_r;
wire main_genericstandalone_crc32_checker_syncfifo_wrport_we;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_wrport_dat_w;
wire main_genericstandalone_crc32_checker_syncfifo_do_read;
wire [2:0] main_genericstandalone_crc32_checker_syncfifo_rdport_adr;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_rdport_dat_r;
wire [7:0] main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_data;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_last_be;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_error;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_in_eop;
wire [7:0] main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_data;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_last_be;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_error;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_out_eop;
reg main_genericstandalone_crc32_checker_fifo_reset;
wire main_genericstandalone_crc32_checker_fifo_in;
wire main_genericstandalone_crc32_checker_fifo_out;
wire main_genericstandalone_crc32_checker_fifo_full;
wire main_genericstandalone_ps_preamble_error_i;
wire main_genericstandalone_ps_preamble_error_o;
reg main_genericstandalone_ps_preamble_error_toggle_i = 1'd0;
wire main_genericstandalone_ps_preamble_error_toggle_o;
reg main_genericstandalone_ps_preamble_error_toggle_o_r = 1'd0;
wire main_genericstandalone_ps_crc_error_i;
wire main_genericstandalone_ps_crc_error_o;
reg main_genericstandalone_ps_crc_error_toggle_i = 1'd0;
wire main_genericstandalone_ps_crc_error_toggle_o;
reg main_genericstandalone_ps_crc_error_toggle_o_r = 1'd0;
wire main_genericstandalone_padding_inserter_sink_stb;
reg main_genericstandalone_padding_inserter_sink_ack;
wire main_genericstandalone_padding_inserter_sink_last;
wire main_genericstandalone_padding_inserter_sink_eop;
wire [7:0] main_genericstandalone_padding_inserter_sink_payload_data;
wire main_genericstandalone_padding_inserter_sink_payload_last_be;
wire main_genericstandalone_padding_inserter_sink_payload_error;
reg main_genericstandalone_padding_inserter_source_stb;
wire main_genericstandalone_padding_inserter_source_ack;
reg main_genericstandalone_padding_inserter_source_last;
reg main_genericstandalone_padding_inserter_source_eop;
reg [7:0] main_genericstandalone_padding_inserter_source_payload_data;
reg main_genericstandalone_padding_inserter_source_payload_last_be;
reg main_genericstandalone_padding_inserter_source_payload_error;
reg [15:0] main_genericstandalone_padding_inserter_counter = 16'd1;
wire main_genericstandalone_padding_inserter_counter_done;
reg main_genericstandalone_padding_inserter_counter_reset;
reg main_genericstandalone_padding_inserter_counter_ce;
wire main_genericstandalone_padding_checker_sink_stb;
wire main_genericstandalone_padding_checker_sink_ack;
wire main_genericstandalone_padding_checker_sink_last;
wire main_genericstandalone_padding_checker_sink_eop;
wire [7:0] main_genericstandalone_padding_checker_sink_payload_data;
wire main_genericstandalone_padding_checker_sink_payload_last_be;
wire main_genericstandalone_padding_checker_sink_payload_error;
wire main_genericstandalone_padding_checker_source_stb;
wire main_genericstandalone_padding_checker_source_ack;
wire main_genericstandalone_padding_checker_source_last;
wire main_genericstandalone_padding_checker_source_eop;
wire [7:0] main_genericstandalone_padding_checker_source_payload_data;
wire main_genericstandalone_padding_checker_source_payload_last_be;
wire main_genericstandalone_padding_checker_source_payload_error;
wire main_genericstandalone_tx_last_be_sink_stb;
wire main_genericstandalone_tx_last_be_sink_ack;
wire main_genericstandalone_tx_last_be_sink_last;
wire main_genericstandalone_tx_last_be_sink_eop;
wire [7:0] main_genericstandalone_tx_last_be_sink_payload_data;
wire main_genericstandalone_tx_last_be_sink_payload_last_be;
wire main_genericstandalone_tx_last_be_sink_payload_error;
wire main_genericstandalone_tx_last_be_source_stb;
wire main_genericstandalone_tx_last_be_source_ack;
reg main_genericstandalone_tx_last_be_source_last = 1'd0;
wire main_genericstandalone_tx_last_be_source_eop;
wire [7:0] main_genericstandalone_tx_last_be_source_payload_data;
reg main_genericstandalone_tx_last_be_source_payload_last_be = 1'd0;
reg main_genericstandalone_tx_last_be_source_payload_error = 1'd0;
reg main_genericstandalone_tx_last_be_ongoing = 1'd1;
wire main_genericstandalone_rx_last_be_sink_stb;
wire main_genericstandalone_rx_last_be_sink_ack;
wire main_genericstandalone_rx_last_be_sink_last;
wire main_genericstandalone_rx_last_be_sink_eop;
wire [7:0] main_genericstandalone_rx_last_be_sink_payload_data;
wire main_genericstandalone_rx_last_be_sink_payload_last_be;
wire main_genericstandalone_rx_last_be_sink_payload_error;
wire main_genericstandalone_rx_last_be_source_stb;
wire main_genericstandalone_rx_last_be_source_ack;
wire main_genericstandalone_rx_last_be_source_last;
wire main_genericstandalone_rx_last_be_source_eop;
wire [7:0] main_genericstandalone_rx_last_be_source_payload_data;
reg main_genericstandalone_rx_last_be_source_payload_last_be;
wire main_genericstandalone_rx_last_be_source_payload_error;
wire main_genericstandalone_tx_converter_sink_sink_stb;
wire main_genericstandalone_tx_converter_sink_sink_ack;
wire main_genericstandalone_tx_converter_sink_sink_last;
wire main_genericstandalone_tx_converter_sink_sink_eop;
wire [63:0] main_genericstandalone_tx_converter_sink_sink_payload_data;
wire [7:0] main_genericstandalone_tx_converter_sink_sink_payload_last_be;
wire [7:0] main_genericstandalone_tx_converter_sink_sink_payload_error;
wire main_genericstandalone_tx_converter_source_source_stb;
wire main_genericstandalone_tx_converter_source_source_ack;
wire main_genericstandalone_tx_converter_source_source_last;
wire main_genericstandalone_tx_converter_source_source_eop;
wire [7:0] main_genericstandalone_tx_converter_source_source_payload_data;
wire main_genericstandalone_tx_converter_source_source_payload_last_be;
wire main_genericstandalone_tx_converter_source_source_payload_error;
wire main_genericstandalone_tx_converter_converter_sink_stb;
wire main_genericstandalone_tx_converter_converter_sink_ack;
wire main_genericstandalone_tx_converter_converter_sink_last;
wire main_genericstandalone_tx_converter_converter_sink_eop;
reg [79:0] main_genericstandalone_tx_converter_converter_sink_payload_data;
wire main_genericstandalone_tx_converter_converter_source_stb;
wire main_genericstandalone_tx_converter_converter_source_ack;
wire main_genericstandalone_tx_converter_converter_source_last;
wire main_genericstandalone_tx_converter_converter_source_eop;
reg [9:0] main_genericstandalone_tx_converter_converter_source_payload_data;
reg [2:0] main_genericstandalone_tx_converter_converter_mux = 3'd0;
wire main_genericstandalone_tx_converter_converter_last;
wire main_genericstandalone_rx_converter_sink_sink_stb;
wire main_genericstandalone_rx_converter_sink_sink_ack;
wire main_genericstandalone_rx_converter_sink_sink_last;
wire main_genericstandalone_rx_converter_sink_sink_eop;
wire [7:0] main_genericstandalone_rx_converter_sink_sink_payload_data;
wire main_genericstandalone_rx_converter_sink_sink_payload_last_be;
wire main_genericstandalone_rx_converter_sink_sink_payload_error;
wire main_genericstandalone_rx_converter_source_source_stb;
wire main_genericstandalone_rx_converter_source_source_ack;
wire main_genericstandalone_rx_converter_source_source_last;
wire main_genericstandalone_rx_converter_source_source_eop;
reg [63:0] main_genericstandalone_rx_converter_source_source_payload_data;
reg [7:0] main_genericstandalone_rx_converter_source_source_payload_last_be;
reg [7:0] main_genericstandalone_rx_converter_source_source_payload_error;
wire main_genericstandalone_rx_converter_converter_sink_stb;
wire main_genericstandalone_rx_converter_converter_sink_ack;
wire main_genericstandalone_rx_converter_converter_sink_last;
wire main_genericstandalone_rx_converter_converter_sink_eop;
wire [9:0] main_genericstandalone_rx_converter_converter_sink_payload_data;
wire main_genericstandalone_rx_converter_converter_source_stb;
wire main_genericstandalone_rx_converter_converter_source_ack;
wire main_genericstandalone_rx_converter_converter_source_last;
reg main_genericstandalone_rx_converter_converter_source_eop = 1'd0;
reg [79:0] main_genericstandalone_rx_converter_converter_source_payload_data = 80'd0;
reg [2:0] main_genericstandalone_rx_converter_converter_demux = 3'd0;
wire main_genericstandalone_rx_converter_converter_load_part;
reg main_genericstandalone_rx_converter_converter_strobe_all = 1'd0;
wire main_genericstandalone_tx_cdc_sink_stb;
wire main_genericstandalone_tx_cdc_sink_ack;
wire main_genericstandalone_tx_cdc_sink_last;
wire main_genericstandalone_tx_cdc_sink_eop;
wire [63:0] main_genericstandalone_tx_cdc_sink_payload_data;
wire [7:0] main_genericstandalone_tx_cdc_sink_payload_last_be;
wire [7:0] main_genericstandalone_tx_cdc_sink_payload_error;
wire main_genericstandalone_tx_cdc_source_stb;
wire main_genericstandalone_tx_cdc_source_ack;
reg main_genericstandalone_tx_cdc_source_last = 1'd0;
wire main_genericstandalone_tx_cdc_source_eop;
wire [63:0] main_genericstandalone_tx_cdc_source_payload_data;
wire [7:0] main_genericstandalone_tx_cdc_source_payload_last_be;
wire [7:0] main_genericstandalone_tx_cdc_source_payload_error;
wire main_genericstandalone_tx_cdc_asyncfifo_we;
wire main_genericstandalone_tx_cdc_asyncfifo_writable;
wire main_genericstandalone_tx_cdc_asyncfifo_re;
wire main_genericstandalone_tx_cdc_asyncfifo_readable;
wire [80:0] main_genericstandalone_tx_cdc_asyncfifo_din;
wire [80:0] main_genericstandalone_tx_cdc_asyncfifo_dout;
wire main_genericstandalone_tx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] main_genericstandalone_tx_cdc_graycounter0_q = 7'd0;
wire [6:0] main_genericstandalone_tx_cdc_graycounter0_q_next;
reg [6:0] main_genericstandalone_tx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] main_genericstandalone_tx_cdc_graycounter0_q_next_binary;
wire main_genericstandalone_tx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] main_genericstandalone_tx_cdc_graycounter1_q = 7'd0;
wire [6:0] main_genericstandalone_tx_cdc_graycounter1_q_next;
reg [6:0] main_genericstandalone_tx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] main_genericstandalone_tx_cdc_graycounter1_q_next_binary;
wire [6:0] main_genericstandalone_tx_cdc_produce_rdomain;
wire [6:0] main_genericstandalone_tx_cdc_consume_wdomain;
wire [5:0] main_genericstandalone_tx_cdc_wrport_adr;
wire [80:0] main_genericstandalone_tx_cdc_wrport_dat_r;
wire main_genericstandalone_tx_cdc_wrport_we;
wire [80:0] main_genericstandalone_tx_cdc_wrport_dat_w;
wire [5:0] main_genericstandalone_tx_cdc_rdport_adr;
wire [80:0] main_genericstandalone_tx_cdc_rdport_dat_r;
wire [63:0] main_genericstandalone_tx_cdc_fifo_in_payload_data;
wire [7:0] main_genericstandalone_tx_cdc_fifo_in_payload_last_be;
wire [7:0] main_genericstandalone_tx_cdc_fifo_in_payload_error;
wire main_genericstandalone_tx_cdc_fifo_in_eop;
wire [63:0] main_genericstandalone_tx_cdc_fifo_out_payload_data;
wire [7:0] main_genericstandalone_tx_cdc_fifo_out_payload_last_be;
wire [7:0] main_genericstandalone_tx_cdc_fifo_out_payload_error;
wire main_genericstandalone_tx_cdc_fifo_out_eop;
wire main_genericstandalone_rx_cdc_sink_stb;
wire main_genericstandalone_rx_cdc_sink_ack;
wire main_genericstandalone_rx_cdc_sink_last;
wire main_genericstandalone_rx_cdc_sink_eop;
wire [63:0] main_genericstandalone_rx_cdc_sink_payload_data;
wire [7:0] main_genericstandalone_rx_cdc_sink_payload_last_be;
wire [7:0] main_genericstandalone_rx_cdc_sink_payload_error;
wire main_genericstandalone_rx_cdc_source_stb;
wire main_genericstandalone_rx_cdc_source_ack;
reg main_genericstandalone_rx_cdc_source_last = 1'd0;
wire main_genericstandalone_rx_cdc_source_eop;
wire [63:0] main_genericstandalone_rx_cdc_source_payload_data;
wire [7:0] main_genericstandalone_rx_cdc_source_payload_last_be;
wire [7:0] main_genericstandalone_rx_cdc_source_payload_error;
wire main_genericstandalone_rx_cdc_asyncfifo_we;
wire main_genericstandalone_rx_cdc_asyncfifo_writable;
wire main_genericstandalone_rx_cdc_asyncfifo_re;
wire main_genericstandalone_rx_cdc_asyncfifo_readable;
wire [80:0] main_genericstandalone_rx_cdc_asyncfifo_din;
wire [80:0] main_genericstandalone_rx_cdc_asyncfifo_dout;
wire main_genericstandalone_rx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] main_genericstandalone_rx_cdc_graycounter0_q = 7'd0;
wire [6:0] main_genericstandalone_rx_cdc_graycounter0_q_next;
reg [6:0] main_genericstandalone_rx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] main_genericstandalone_rx_cdc_graycounter0_q_next_binary;
wire main_genericstandalone_rx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] main_genericstandalone_rx_cdc_graycounter1_q = 7'd0;
wire [6:0] main_genericstandalone_rx_cdc_graycounter1_q_next;
reg [6:0] main_genericstandalone_rx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] main_genericstandalone_rx_cdc_graycounter1_q_next_binary;
wire [6:0] main_genericstandalone_rx_cdc_produce_rdomain;
wire [6:0] main_genericstandalone_rx_cdc_consume_wdomain;
wire [5:0] main_genericstandalone_rx_cdc_wrport_adr;
wire [80:0] main_genericstandalone_rx_cdc_wrport_dat_r;
wire main_genericstandalone_rx_cdc_wrport_we;
wire [80:0] main_genericstandalone_rx_cdc_wrport_dat_w;
wire [5:0] main_genericstandalone_rx_cdc_rdport_adr;
wire [80:0] main_genericstandalone_rx_cdc_rdport_dat_r;
wire [63:0] main_genericstandalone_rx_cdc_fifo_in_payload_data;
wire [7:0] main_genericstandalone_rx_cdc_fifo_in_payload_last_be;
wire [7:0] main_genericstandalone_rx_cdc_fifo_in_payload_error;
wire main_genericstandalone_rx_cdc_fifo_in_eop;
wire [63:0] main_genericstandalone_rx_cdc_fifo_out_payload_data;
wire [7:0] main_genericstandalone_rx_cdc_fifo_out_payload_last_be;
wire [7:0] main_genericstandalone_rx_cdc_fifo_out_payload_error;
wire main_genericstandalone_rx_cdc_fifo_out_eop;
wire main_genericstandalone_sink_sink_stb;
wire main_genericstandalone_sink_sink_ack;
wire main_genericstandalone_sink_sink_last;
wire main_genericstandalone_sink_sink_eop;
wire [63:0] main_genericstandalone_sink_sink_payload_data;
wire [7:0] main_genericstandalone_sink_sink_payload_last_be;
wire [7:0] main_genericstandalone_sink_sink_payload_error;
wire main_genericstandalone_source_source_stb;
wire main_genericstandalone_source_source_ack;
wire main_genericstandalone_source_source_last;
wire main_genericstandalone_source_source_eop;
wire [63:0] main_genericstandalone_source_source_payload_data;
wire [7:0] main_genericstandalone_source_source_payload_last_be;
wire [7:0] main_genericstandalone_source_source_payload_error;
wire [28:0] main_genericstandalone_bus_bus_adr;
wire [63:0] main_genericstandalone_bus_bus_dat_w;
wire [63:0] main_genericstandalone_bus_bus_dat_r;
wire [7:0] main_genericstandalone_bus_bus_sel;
wire main_genericstandalone_bus_bus_cyc;
wire main_genericstandalone_bus_bus_stb;
wire main_genericstandalone_bus_bus_ack;
wire main_genericstandalone_bus_bus_we;
wire [2:0] main_genericstandalone_bus_bus_cti;
wire [1:0] main_genericstandalone_bus_bus_bte;
wire main_genericstandalone_bus_bus_err;
wire main_genericstandalone_sram8_sink_stb;
reg main_genericstandalone_sram9_sink_ack = 1'd1;
wire main_genericstandalone_sram10_sink_last;
wire main_genericstandalone_sram11_sink_eop;
wire [63:0] main_genericstandalone_sram12_sink_payload_data;
wire [7:0] main_genericstandalone_sram13_sink_payload_last_be;
wire [7:0] main_genericstandalone_sram14_sink_payload_error;
wire [1:0] main_genericstandalone_sram15_status;
wire [10:0] main_genericstandalone_sram16_status;
reg [31:0] main_genericstandalone_sram17_status = 32'd0;
wire main_genericstandalone_sram18_irq;
wire main_genericstandalone_sram19_status;
wire main_genericstandalone_sram20_pending;
wire main_genericstandalone_sram21_trigger;
reg main_genericstandalone_sram22_clear;
wire main_genericstandalone_sram23_status_re;
wire main_genericstandalone_sram24_status_r;
wire main_genericstandalone_sram25_status_w;
wire main_genericstandalone_sram26_pending_re;
wire main_genericstandalone_sram27_pending_r;
wire main_genericstandalone_sram28_pending_w;
reg main_genericstandalone_sram29_storage_full = 1'd0;
wire main_genericstandalone_sram30_storage;
reg main_genericstandalone_sram31_re = 1'd0;
reg [3:0] main_genericstandalone_decoded;
reg [10:0] main_genericstandalone_sram33_counter = 11'd0;
reg main_genericstandalone_sram34_counter_reset;
reg main_genericstandalone_sram35_counter_ce;
reg [1:0] main_genericstandalone_slot = 2'd0;
reg main_genericstandalone_slot_ce;
reg main_genericstandalone_ongoing;
reg main_genericstandalone_sram39_sink_stb;
wire main_genericstandalone_sram40_sink_ack;
reg main_genericstandalone_sram41_sink_eop = 1'd0;
wire [1:0] main_genericstandalone_sram42_sink_payload_slot;
wire [10:0] main_genericstandalone_sram43_sink_payload_length;
wire main_genericstandalone_sram44_source_stb;
wire main_genericstandalone_sram45_source_ack;
wire main_genericstandalone_sram46_source_eop;
wire [1:0] main_genericstandalone_sram47_source_payload_slot;
wire [10:0] main_genericstandalone_sram48_source_payload_length;
wire main_genericstandalone_sram49_we;
wire main_genericstandalone_sram50_writable;
wire main_genericstandalone_sram51_re;
wire main_genericstandalone_sram52_readable;
wire [13:0] main_genericstandalone_sram53_din;
wire [13:0] main_genericstandalone_sram54_dout;
reg [2:0] main_genericstandalone_sram55_level = 3'd0;
reg main_genericstandalone_sram56_replace = 1'd0;
reg [1:0] main_genericstandalone_sram57_produce = 2'd0;
reg [1:0] main_genericstandalone_sram58_consume = 2'd0;
reg [1:0] main_genericstandalone_sram59_adr;
wire [13:0] main_genericstandalone_sram60_dat_r;
wire main_genericstandalone_sram61_we;
wire [13:0] main_genericstandalone_sram62_dat_w;
wire main_genericstandalone_sram63_do_read;
wire [1:0] main_genericstandalone_sram64_adr;
wire [13:0] main_genericstandalone_sram65_dat_r;
wire [1:0] main_genericstandalone_sram66_fifo_in_payload_slot;
wire [10:0] main_genericstandalone_sram67_fifo_in_payload_length;
wire main_genericstandalone_sram68_fifo_in_eop;
wire [1:0] main_genericstandalone_sram69_fifo_out_payload_slot;
wire [10:0] main_genericstandalone_sram70_fifo_out_payload_length;
wire main_genericstandalone_sram71_fifo_out_eop;
reg [7:0] main_genericstandalone_sram72_adr;
wire [63:0] main_genericstandalone_sram73_dat_r;
reg main_genericstandalone_sram74_we;
reg [63:0] main_genericstandalone_sram75_dat_w;
reg [7:0] main_genericstandalone_sram76_adr;
wire [63:0] main_genericstandalone_sram77_dat_r;
reg main_genericstandalone_sram78_we;
reg [63:0] main_genericstandalone_sram79_dat_w;
reg [7:0] main_genericstandalone_sram80_adr;
wire [63:0] main_genericstandalone_sram81_dat_r;
reg main_genericstandalone_sram82_we;
reg [63:0] main_genericstandalone_sram83_dat_w;
reg [7:0] main_genericstandalone_sram84_adr;
wire [63:0] main_genericstandalone_sram85_dat_r;
reg main_genericstandalone_sram86_we;
reg [63:0] main_genericstandalone_sram87_dat_w;
reg main_genericstandalone_sram88_source_stb;
wire main_genericstandalone_sram89_source_ack;
reg main_genericstandalone_sram90_source_last = 1'd0;
reg main_genericstandalone_sram91_source_eop;
reg [63:0] main_genericstandalone_sram92_source_payload_data;
reg [7:0] main_genericstandalone_sram93_source_payload_last_be;
reg [7:0] main_genericstandalone_sram94_source_payload_error = 8'd0;
wire main_genericstandalone_start_re;
wire main_genericstandalone_start_r;
reg main_genericstandalone_start_w = 1'd0;
wire main_genericstandalone_sram98_status;
reg [1:0] main_genericstandalone_sram99_storage_full = 2'd0;
wire [1:0] main_genericstandalone_sram100_storage;
reg main_genericstandalone_sram101_re = 1'd0;
reg [10:0] main_genericstandalone_sram102_storage_full = 11'd0;
wire [10:0] main_genericstandalone_sram103_storage;
reg main_genericstandalone_sram104_re = 1'd0;
wire main_genericstandalone_sram105_irq;
wire main_genericstandalone_sram106_status;
reg main_genericstandalone_sram107_pending = 1'd0;
reg main_genericstandalone_sram108_trigger;
reg main_genericstandalone_sram109_clear;
wire main_genericstandalone_sram110_status_re;
wire main_genericstandalone_sram111_status_r;
wire main_genericstandalone_sram112_status_w;
wire main_genericstandalone_sram113_pending_re;
wire main_genericstandalone_sram114_pending_r;
wire main_genericstandalone_sram115_pending_w;
reg main_genericstandalone_sram116_storage_full = 1'd0;
wire main_genericstandalone_sram117_storage;
reg main_genericstandalone_sram118_re = 1'd0;
wire main_genericstandalone_sram119_sink_stb;
wire main_genericstandalone_sram120_sink_ack;
reg main_genericstandalone_sram121_sink_eop = 1'd0;
wire [1:0] main_genericstandalone_sram122_sink_payload_slot;
wire [10:0] main_genericstandalone_sram123_sink_payload_length;
wire main_genericstandalone_sram124_source_stb;
reg main_genericstandalone_sram125_source_ack;
wire main_genericstandalone_sram126_source_eop;
wire [1:0] main_genericstandalone_sram127_source_payload_slot;
wire [10:0] main_genericstandalone_sram128_source_payload_length;
wire main_genericstandalone_sram129_we;
wire main_genericstandalone_sram130_writable;
wire main_genericstandalone_sram131_re;
wire main_genericstandalone_sram132_readable;
wire [13:0] main_genericstandalone_sram133_din;
wire [13:0] main_genericstandalone_sram134_dout;
reg [2:0] main_genericstandalone_sram135_level = 3'd0;
reg main_genericstandalone_sram136_replace = 1'd0;
reg [1:0] main_genericstandalone_sram137_produce = 2'd0;
reg [1:0] main_genericstandalone_sram138_consume = 2'd0;
reg [1:0] main_genericstandalone_sram139_adr;
wire [13:0] main_genericstandalone_sram140_dat_r;
wire main_genericstandalone_sram141_we;
wire [13:0] main_genericstandalone_sram142_dat_w;
wire main_genericstandalone_sram143_do_read;
wire [1:0] main_genericstandalone_sram144_adr;
wire [13:0] main_genericstandalone_sram145_dat_r;
wire [1:0] main_genericstandalone_sram146_fifo_in_payload_slot;
wire [10:0] main_genericstandalone_sram147_fifo_in_payload_length;
wire main_genericstandalone_sram148_fifo_in_eop;
wire [1:0] main_genericstandalone_sram149_fifo_out_payload_slot;
wire [10:0] main_genericstandalone_sram150_fifo_out_payload_length;
wire main_genericstandalone_sram151_fifo_out_eop;
reg [10:0] main_genericstandalone_sram152_counter = 11'd0;
reg main_genericstandalone_sram153_counter_reset;
reg main_genericstandalone_sram154_counter_ce;
wire main_genericstandalone_last;
reg main_genericstandalone_last_d = 1'd0;
reg [7:0] main_genericstandalone_encoded;
wire [7:0] main_genericstandalone_sram158_adr;
wire [63:0] main_genericstandalone_sram159_dat_r;
wire [7:0] main_genericstandalone_sram160_adr;
wire [63:0] main_genericstandalone_sram161_dat_r;
wire [7:0] main_genericstandalone_sram162_adr;
wire [63:0] main_genericstandalone_sram163_dat_r;
wire [7:0] main_genericstandalone_sram164_adr;
wire [63:0] main_genericstandalone_sram165_dat_r;
wire main_genericstandalone_sram166_irq;
wire [28:0] main_genericstandalone_sram0_bus_adr;
wire [63:0] main_genericstandalone_sram0_bus_dat_w;
wire [63:0] main_genericstandalone_sram0_bus_dat_r;
wire [7:0] main_genericstandalone_sram0_bus_sel;
wire main_genericstandalone_sram0_bus_cyc;
wire main_genericstandalone_sram0_bus_stb;
reg main_genericstandalone_sram0_bus_ack = 1'd0;
wire main_genericstandalone_sram0_bus_we;
wire [2:0] main_genericstandalone_sram0_bus_cti;
wire [1:0] main_genericstandalone_sram0_bus_bte;
reg main_genericstandalone_sram0_bus_err = 1'd0;
wire [7:0] main_genericstandalone_sram0_adr;
wire [63:0] main_genericstandalone_sram0_dat_r;
wire [28:0] main_genericstandalone_sram1_bus_adr;
wire [63:0] main_genericstandalone_sram1_bus_dat_w;
wire [63:0] main_genericstandalone_sram1_bus_dat_r;
wire [7:0] main_genericstandalone_sram1_bus_sel;
wire main_genericstandalone_sram1_bus_cyc;
wire main_genericstandalone_sram1_bus_stb;
reg main_genericstandalone_sram1_bus_ack = 1'd0;
wire main_genericstandalone_sram1_bus_we;
wire [2:0] main_genericstandalone_sram1_bus_cti;
wire [1:0] main_genericstandalone_sram1_bus_bte;
reg main_genericstandalone_sram1_bus_err = 1'd0;
wire [7:0] main_genericstandalone_sram1_adr;
wire [63:0] main_genericstandalone_sram1_dat_r;
wire [28:0] main_genericstandalone_sram2_bus_adr;
wire [63:0] main_genericstandalone_sram2_bus_dat_w;
wire [63:0] main_genericstandalone_sram2_bus_dat_r;
wire [7:0] main_genericstandalone_sram2_bus_sel;
wire main_genericstandalone_sram2_bus_cyc;
wire main_genericstandalone_sram2_bus_stb;
reg main_genericstandalone_sram2_bus_ack = 1'd0;
wire main_genericstandalone_sram2_bus_we;
wire [2:0] main_genericstandalone_sram2_bus_cti;
wire [1:0] main_genericstandalone_sram2_bus_bte;
reg main_genericstandalone_sram2_bus_err = 1'd0;
wire [7:0] main_genericstandalone_sram2_adr;
wire [63:0] main_genericstandalone_sram2_dat_r;
wire [28:0] main_genericstandalone_sram3_bus_adr;
wire [63:0] main_genericstandalone_sram3_bus_dat_w;
wire [63:0] main_genericstandalone_sram3_bus_dat_r;
wire [7:0] main_genericstandalone_sram3_bus_sel;
wire main_genericstandalone_sram3_bus_cyc;
wire main_genericstandalone_sram3_bus_stb;
reg main_genericstandalone_sram3_bus_ack = 1'd0;
wire main_genericstandalone_sram3_bus_we;
wire [2:0] main_genericstandalone_sram3_bus_cti;
wire [1:0] main_genericstandalone_sram3_bus_bte;
reg main_genericstandalone_sram3_bus_err = 1'd0;
wire [7:0] main_genericstandalone_sram3_adr;
wire [63:0] main_genericstandalone_sram3_dat_r;
wire [28:0] main_genericstandalone_sram4_bus_adr;
wire [63:0] main_genericstandalone_sram4_bus_dat_w;
wire [63:0] main_genericstandalone_sram4_bus_dat_r;
wire [7:0] main_genericstandalone_sram4_bus_sel;
wire main_genericstandalone_sram4_bus_cyc;
wire main_genericstandalone_sram4_bus_stb;
reg main_genericstandalone_sram4_bus_ack = 1'd0;
wire main_genericstandalone_sram4_bus_we;
wire [2:0] main_genericstandalone_sram4_bus_cti;
wire [1:0] main_genericstandalone_sram4_bus_bte;
reg main_genericstandalone_sram4_bus_err = 1'd0;
wire [7:0] main_genericstandalone_sram4_adr;
wire [63:0] main_genericstandalone_sram4_dat_r;
reg [7:0] main_genericstandalone_sram4_we;
wire [63:0] main_genericstandalone_sram4_dat_w;
wire [28:0] main_genericstandalone_sram5_bus_adr;
wire [63:0] main_genericstandalone_sram5_bus_dat_w;
wire [63:0] main_genericstandalone_sram5_bus_dat_r;
wire [7:0] main_genericstandalone_sram5_bus_sel;
wire main_genericstandalone_sram5_bus_cyc;
wire main_genericstandalone_sram5_bus_stb;
reg main_genericstandalone_sram5_bus_ack = 1'd0;
wire main_genericstandalone_sram5_bus_we;
wire [2:0] main_genericstandalone_sram5_bus_cti;
wire [1:0] main_genericstandalone_sram5_bus_bte;
reg main_genericstandalone_sram5_bus_err = 1'd0;
wire [7:0] main_genericstandalone_sram5_adr;
wire [63:0] main_genericstandalone_sram5_dat_r;
reg [7:0] main_genericstandalone_sram5_we;
wire [63:0] main_genericstandalone_sram5_dat_w;
wire [28:0] main_genericstandalone_sram6_bus_adr;
wire [63:0] main_genericstandalone_sram6_bus_dat_w;
wire [63:0] main_genericstandalone_sram6_bus_dat_r;
wire [7:0] main_genericstandalone_sram6_bus_sel;
wire main_genericstandalone_sram6_bus_cyc;
wire main_genericstandalone_sram6_bus_stb;
reg main_genericstandalone_sram6_bus_ack = 1'd0;
wire main_genericstandalone_sram6_bus_we;
wire [2:0] main_genericstandalone_sram6_bus_cti;
wire [1:0] main_genericstandalone_sram6_bus_bte;
reg main_genericstandalone_sram6_bus_err = 1'd0;
wire [7:0] main_genericstandalone_sram6_adr;
wire [63:0] main_genericstandalone_sram6_dat_r;
reg [7:0] main_genericstandalone_sram6_we;
wire [63:0] main_genericstandalone_sram6_dat_w;
wire [28:0] main_genericstandalone_sram7_bus_adr;
wire [63:0] main_genericstandalone_sram7_bus_dat_w;
wire [63:0] main_genericstandalone_sram7_bus_dat_r;
wire [7:0] main_genericstandalone_sram7_bus_sel;
wire main_genericstandalone_sram7_bus_cyc;
wire main_genericstandalone_sram7_bus_stb;
reg main_genericstandalone_sram7_bus_ack = 1'd0;
wire main_genericstandalone_sram7_bus_we;
wire [2:0] main_genericstandalone_sram7_bus_cti;
wire [1:0] main_genericstandalone_sram7_bus_bte;
reg main_genericstandalone_sram7_bus_err = 1'd0;
wire [7:0] main_genericstandalone_sram7_adr;
wire [63:0] main_genericstandalone_sram7_dat_r;
reg [7:0] main_genericstandalone_sram7_we;
wire [63:0] main_genericstandalone_sram7_dat_w;
reg [7:0] main_genericstandalone_slave_sel;
reg [7:0] main_genericstandalone_slave_sel_r = 8'd0;
reg main_genericstandalone_kernel_cpu_storage_full = 1'd1;
wire main_genericstandalone_kernel_cpu_storage;
reg main_genericstandalone_kernel_cpu_re = 1'd0;
wire sys_kernel_clk;
wire sys_kernel_rst;
wire [28:0] main_genericstandalone_kernel_cpu_ibus_adr;
wire [63:0] main_genericstandalone_kernel_cpu_ibus_dat_w;
wire [63:0] main_genericstandalone_kernel_cpu_ibus_dat_r;
wire [7:0] main_genericstandalone_kernel_cpu_ibus_sel;
wire main_genericstandalone_kernel_cpu_ibus_cyc;
wire main_genericstandalone_kernel_cpu_ibus_stb;
wire main_genericstandalone_kernel_cpu_ibus_ack;
wire main_genericstandalone_kernel_cpu_ibus_we;
wire [2:0] main_genericstandalone_kernel_cpu_ibus_cti;
wire [1:0] main_genericstandalone_kernel_cpu_ibus_bte;
wire main_genericstandalone_kernel_cpu_ibus_err;
wire [28:0] main_genericstandalone_kernel_cpu_dbus_adr;
wire [63:0] main_genericstandalone_kernel_cpu_dbus_dat_w;
wire [63:0] main_genericstandalone_kernel_cpu_dbus_dat_r;
wire [7:0] main_genericstandalone_kernel_cpu_dbus_sel;
wire main_genericstandalone_kernel_cpu_dbus_cyc;
wire main_genericstandalone_kernel_cpu_dbus_stb;
wire main_genericstandalone_kernel_cpu_dbus_ack;
wire main_genericstandalone_kernel_cpu_dbus_we;
wire [2:0] main_genericstandalone_kernel_cpu_dbus_cti;
wire [1:0] main_genericstandalone_kernel_cpu_dbus_bte;
wire main_genericstandalone_kernel_cpu_dbus_err;
reg [31:0] main_genericstandalone_kernel_cpu_interrupt = 32'd0;
wire [28:0] main_genericstandalone_kernel_cpu_wb_sdram_adr;
wire [63:0] main_genericstandalone_kernel_cpu_wb_sdram_dat_w;
wire [63:0] main_genericstandalone_kernel_cpu_wb_sdram_dat_r;
wire [7:0] main_genericstandalone_kernel_cpu_wb_sdram_sel;
wire main_genericstandalone_kernel_cpu_wb_sdram_cyc;
wire main_genericstandalone_kernel_cpu_wb_sdram_stb;
wire main_genericstandalone_kernel_cpu_wb_sdram_ack;
wire main_genericstandalone_kernel_cpu_wb_sdram_we;
wire [2:0] main_genericstandalone_kernel_cpu_wb_sdram_cti;
wire [1:0] main_genericstandalone_kernel_cpu_wb_sdram_bte;
wire main_genericstandalone_kernel_cpu_wb_sdram_err;
wire [28:0] main_genericstandalone_mailbox_i1_adr;
wire [31:0] main_genericstandalone_mailbox_i1_dat_w;
reg [31:0] main_genericstandalone_mailbox_i1_dat_r = 32'd0;
wire [3:0] main_genericstandalone_mailbox_i1_sel;
wire main_genericstandalone_mailbox_i1_cyc;
wire main_genericstandalone_mailbox_i1_stb;
reg main_genericstandalone_mailbox_i1_ack = 1'd0;
wire main_genericstandalone_mailbox_i1_we;
wire [2:0] main_genericstandalone_mailbox_i1_cti;
wire [1:0] main_genericstandalone_mailbox_i1_bte;
reg main_genericstandalone_mailbox_i1_err = 1'd0;
wire [28:0] main_genericstandalone_mailbox_i2_adr;
wire [31:0] main_genericstandalone_mailbox_i2_dat_w;
reg [31:0] main_genericstandalone_mailbox_i2_dat_r = 32'd0;
wire [3:0] main_genericstandalone_mailbox_i2_sel;
wire main_genericstandalone_mailbox_i2_cyc;
wire main_genericstandalone_mailbox_i2_stb;
reg main_genericstandalone_mailbox_i2_ack = 1'd0;
wire main_genericstandalone_mailbox_i2_we;
wire [2:0] main_genericstandalone_mailbox_i2_cti;
wire [1:0] main_genericstandalone_mailbox_i2_bte;
reg main_genericstandalone_mailbox_i2_err = 1'd0;
reg [31:0] main_genericstandalone_mailbox0 = 32'd0;
reg [31:0] main_genericstandalone_mailbox1 = 32'd0;
reg [31:0] main_genericstandalone_mailbox2 = 32'd0;
reg [7:0] main_genericstandalone_add_identifier_storage_full = 8'd0;
wire [7:0] main_genericstandalone_add_identifier_storage;
reg main_genericstandalone_add_identifier_re = 1'd0;
wire [7:0] main_genericstandalone_add_identifier_status;
reg main_genericstandalone_error_led_storage_full = 1'd0;
wire main_genericstandalone_error_led_storage;
reg main_genericstandalone_error_led_re = 1'd0;
wire main_genericstandalone_cdr_clk;
wire main_genericstandalone_cdr_clk_buf;
wire main_genericstandalone_rtiosyscrg_mmcm_fb_in;
wire main_genericstandalone_rtiosyscrg_mmcm_fb_out;
wire main_genericstandalone_rtiosyscrg_mmcm_locked;
wire main_genericstandalone_rtiosyscrg_mmcm_sys;
wire main_genericstandalone_rtiosyscrg_mmcm_sys4x;
wire main_genericstandalone_rtiosyscrg_mmcm_sys4x_dqs;
wire main_genericstandalone_rtiosyscrg_async_reset;
wire main_genericstandalone_rtiosyscrg_rst_meta;
wire main_genericstandalone_rtiosyscrg_rst_unbuf;
reg main_genericstandalone_rtiosyscrg_storage_full = 1'd0;
wire main_genericstandalone_rtiosyscrg_storage;
reg main_genericstandalone_rtiosyscrg_re = 1'd0;
wire main_genericstandalone_sma_clkin_se;
wire main_genericstandalone_sma_clkin_buffered;
wire main_genericstandalone_cdr_clk_se;
reg [1:0] main_genericstandalone_i2c_status0;
reg [1:0] main_genericstandalone_i2c_out_storage_full = 2'd0;
wire [1:0] main_genericstandalone_i2c_out_storage;
reg main_genericstandalone_i2c_out_re = 1'd0;
reg [1:0] main_genericstandalone_i2c_oe_storage_full = 2'd0;
wire [1:0] main_genericstandalone_i2c_oe_storage;
reg main_genericstandalone_i2c_oe_re = 1'd0;
wire main_genericstandalone_i2c_tstriple0_o;
wire main_genericstandalone_i2c_tstriple0_oe;
wire main_genericstandalone_i2c_tstriple0_i;
wire main_genericstandalone_i2c_status1;
wire main_genericstandalone_i2c_tstriple1_o;
wire main_genericstandalone_i2c_tstriple1_oe;
wire main_genericstandalone_i2c_tstriple1_i;
wire main_genericstandalone_i2c_status2;
reg [7:0] main_inout_8x0_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x0_serdes_i0;
wire main_inout_8x0_serdes_oe;
wire main_inout_8x0_serdes_ser_in;
wire [7:0] main_inout_8x0_serdes_i1;
wire main_inout_8x0_serdes_ser_out;
wire [7:0] main_inout_8x0_serdes_o1;
wire main_inout_8x0_serdes_t_in;
wire main_inout_8x0_serdes_t_out;
reg main_inout_8x0_inout_8x0_ointerface0_stb = 1'd0;
reg main_inout_8x0_inout_8x0_ointerface0_busy = 1'd0;
reg [1:0] main_inout_8x0_inout_8x0_ointerface0_data = 2'd0;
reg [1:0] main_inout_8x0_inout_8x0_ointerface0_address = 2'd0;
reg [2:0] main_inout_8x0_inout_8x0_ointerface0_fine_ts = 3'd0;
reg main_inout_8x0_inout_8x0_iinterface0_stb = 1'd0;
reg main_inout_8x0_inout_8x0_iinterface0_data = 1'd0;
reg [2:0] main_inout_8x0_inout_8x0_iinterface0_fine_ts = 3'd0;
wire main_inout_8x0_inout_8x0_override_en;
wire main_inout_8x0_inout_8x0_override_o;
wire main_inout_8x0_inout_8x0_override_oe;
(* dont_touch = "true" *) reg main_inout_8x0_inout_8x0_oe = 1'd0;
wire main_inout_8x0_inout_8x0_input_state;
reg main_inout_8x0_inout_8x0_previous_data = 1'd0;
reg main_inout_8x0_inout_8x0_oe_k = 1'd0;
reg [1:0] main_inout_8x0_inout_8x0_sensitivity = 2'd0;
reg main_inout_8x0_inout_8x0_sample = 1'd0;
reg main_inout_8x0_inout_8x0_i_d = 1'd0;
wire [7:0] main_inout_8x0_inout_8x0_i;
reg [2:0] main_inout_8x0_inout_8x0_o;
wire main_inout_8x0_inout_8x0_n;
reg [7:0] main_inout_8x1_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x1_serdes_i0;
wire main_inout_8x1_serdes_oe;
wire main_inout_8x1_serdes_ser_in;
wire [7:0] main_inout_8x1_serdes_i1;
wire main_inout_8x1_serdes_ser_out;
wire [7:0] main_inout_8x1_serdes_o1;
wire main_inout_8x1_serdes_t_in;
wire main_inout_8x1_serdes_t_out;
reg main_inout_8x1_inout_8x1_ointerface1_stb = 1'd0;
reg main_inout_8x1_inout_8x1_ointerface1_busy = 1'd0;
reg [1:0] main_inout_8x1_inout_8x1_ointerface1_data = 2'd0;
reg [1:0] main_inout_8x1_inout_8x1_ointerface1_address = 2'd0;
reg [2:0] main_inout_8x1_inout_8x1_ointerface1_fine_ts = 3'd0;
reg main_inout_8x1_inout_8x1_iinterface1_stb = 1'd0;
reg main_inout_8x1_inout_8x1_iinterface1_data = 1'd0;
reg [2:0] main_inout_8x1_inout_8x1_iinterface1_fine_ts = 3'd0;
wire main_inout_8x1_inout_8x1_override_en;
wire main_inout_8x1_inout_8x1_override_o;
wire main_inout_8x1_inout_8x1_override_oe;
(* dont_touch = "true" *) reg main_inout_8x1_inout_8x1_oe = 1'd0;
wire main_inout_8x1_inout_8x1_input_state;
reg main_inout_8x1_inout_8x1_previous_data = 1'd0;
reg main_inout_8x1_inout_8x1_oe_k = 1'd0;
reg [1:0] main_inout_8x1_inout_8x1_sensitivity = 2'd0;
reg main_inout_8x1_inout_8x1_sample = 1'd0;
reg main_inout_8x1_inout_8x1_i_d = 1'd0;
wire [7:0] main_inout_8x1_inout_8x1_i;
reg [2:0] main_inout_8x1_inout_8x1_o;
wire main_inout_8x1_inout_8x1_n;
reg [7:0] main_inout_8x2_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x2_serdes_i0;
wire main_inout_8x2_serdes_oe;
wire main_inout_8x2_serdes_ser_in;
wire [7:0] main_inout_8x2_serdes_i1;
wire main_inout_8x2_serdes_ser_out;
wire [7:0] main_inout_8x2_serdes_o1;
wire main_inout_8x2_serdes_t_in;
wire main_inout_8x2_serdes_t_out;
reg main_inout_8x2_inout_8x2_ointerface2_stb = 1'd0;
reg main_inout_8x2_inout_8x2_ointerface2_busy = 1'd0;
reg [1:0] main_inout_8x2_inout_8x2_ointerface2_data = 2'd0;
reg [1:0] main_inout_8x2_inout_8x2_ointerface2_address = 2'd0;
reg [2:0] main_inout_8x2_inout_8x2_ointerface2_fine_ts = 3'd0;
reg main_inout_8x2_inout_8x2_iinterface2_stb = 1'd0;
reg main_inout_8x2_inout_8x2_iinterface2_data = 1'd0;
reg [2:0] main_inout_8x2_inout_8x2_iinterface2_fine_ts = 3'd0;
wire main_inout_8x2_inout_8x2_override_en;
wire main_inout_8x2_inout_8x2_override_o;
wire main_inout_8x2_inout_8x2_override_oe;
(* dont_touch = "true" *) reg main_inout_8x2_inout_8x2_oe = 1'd0;
wire main_inout_8x2_inout_8x2_input_state;
reg main_inout_8x2_inout_8x2_previous_data = 1'd0;
reg main_inout_8x2_inout_8x2_oe_k = 1'd0;
reg [1:0] main_inout_8x2_inout_8x2_sensitivity = 2'd0;
reg main_inout_8x2_inout_8x2_sample = 1'd0;
reg main_inout_8x2_inout_8x2_i_d = 1'd0;
wire [7:0] main_inout_8x2_inout_8x2_i;
reg [2:0] main_inout_8x2_inout_8x2_o;
wire main_inout_8x2_inout_8x2_n;
reg [7:0] main_inout_8x3_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x3_serdes_i0;
wire main_inout_8x3_serdes_oe;
wire main_inout_8x3_serdes_ser_in;
wire [7:0] main_inout_8x3_serdes_i1;
wire main_inout_8x3_serdes_ser_out;
wire [7:0] main_inout_8x3_serdes_o1;
wire main_inout_8x3_serdes_t_in;
wire main_inout_8x3_serdes_t_out;
reg main_inout_8x3_inout_8x3_ointerface3_stb = 1'd0;
reg main_inout_8x3_inout_8x3_ointerface3_busy = 1'd0;
reg [1:0] main_inout_8x3_inout_8x3_ointerface3_data = 2'd0;
reg [1:0] main_inout_8x3_inout_8x3_ointerface3_address = 2'd0;
reg [2:0] main_inout_8x3_inout_8x3_ointerface3_fine_ts = 3'd0;
reg main_inout_8x3_inout_8x3_iinterface3_stb = 1'd0;
reg main_inout_8x3_inout_8x3_iinterface3_data = 1'd0;
reg [2:0] main_inout_8x3_inout_8x3_iinterface3_fine_ts = 3'd0;
wire main_inout_8x3_inout_8x3_override_en;
wire main_inout_8x3_inout_8x3_override_o;
wire main_inout_8x3_inout_8x3_override_oe;
(* dont_touch = "true" *) reg main_inout_8x3_inout_8x3_oe = 1'd0;
wire main_inout_8x3_inout_8x3_input_state;
reg main_inout_8x3_inout_8x3_previous_data = 1'd0;
reg main_inout_8x3_inout_8x3_oe_k = 1'd0;
reg [1:0] main_inout_8x3_inout_8x3_sensitivity = 2'd0;
reg main_inout_8x3_inout_8x3_sample = 1'd0;
reg main_inout_8x3_inout_8x3_i_d = 1'd0;
wire [7:0] main_inout_8x3_inout_8x3_i;
reg [2:0] main_inout_8x3_inout_8x3_o;
wire main_inout_8x3_inout_8x3_n;
wire main_output_8x0_ser_out0;
reg [7:0] main_output_8x0_o0 = 8'd0;
reg main_output_8x0_t_in0 = 1'd0;
wire main_output_8x0_t_out0;
reg main_output_8x0_stb0 = 1'd0;
reg main_output_8x0_busy0 = 1'd0;
reg main_output_8x0_data0 = 1'd0;
reg [2:0] main_output_8x0_fine_ts0 = 3'd0;
wire main_output_8x0_override_en0;
wire main_output_8x0_override_o0;
reg main_output_8x0_previous_data0 = 1'd0;
wire main_output_8x1_ser_out0;
reg [7:0] main_output_8x1_o0 = 8'd0;
reg main_output_8x1_t_in0 = 1'd0;
wire main_output_8x1_t_out0;
reg main_output_8x1_stb0 = 1'd0;
reg main_output_8x1_busy0 = 1'd0;
reg main_output_8x1_data0 = 1'd0;
reg [2:0] main_output_8x1_fine_ts0 = 3'd0;
wire main_output_8x1_override_en0;
wire main_output_8x1_override_o0;
reg main_output_8x1_previous_data0 = 1'd0;
wire main_output_8x2_ser_out;
reg [7:0] main_output_8x2_o = 8'd0;
reg main_output_8x2_t_in = 1'd0;
wire main_output_8x2_t_out;
reg main_output_8x2_stb = 1'd0;
reg main_output_8x2_busy = 1'd0;
reg main_output_8x2_data = 1'd0;
reg [2:0] main_output_8x2_fine_ts = 3'd0;
wire main_output_8x2_override_en;
wire main_output_8x2_override_o;
reg main_output_8x2_previous_data = 1'd0;
wire main_output_8x3_ser_out;
reg [7:0] main_output_8x3_o = 8'd0;
reg main_output_8x3_t_in = 1'd0;
wire main_output_8x3_t_out;
reg main_output_8x3_stb = 1'd0;
reg main_output_8x3_busy = 1'd0;
reg main_output_8x3_data = 1'd0;
reg [2:0] main_output_8x3_fine_ts = 3'd0;
wire main_output_8x3_override_en;
wire main_output_8x3_override_o;
reg main_output_8x3_previous_data = 1'd0;
wire main_output_8x4_ser_out;
reg [7:0] main_output_8x4_o = 8'd0;
reg main_output_8x4_t_in = 1'd0;
wire main_output_8x4_t_out;
reg main_output_8x4_stb = 1'd0;
reg main_output_8x4_busy = 1'd0;
reg main_output_8x4_data = 1'd0;
reg [2:0] main_output_8x4_fine_ts = 3'd0;
wire main_output_8x4_override_en;
wire main_output_8x4_override_o;
reg main_output_8x4_previous_data = 1'd0;
wire main_output_8x5_ser_out;
reg [7:0] main_output_8x5_o = 8'd0;
reg main_output_8x5_t_in = 1'd0;
wire main_output_8x5_t_out;
reg main_output_8x5_stb = 1'd0;
reg main_output_8x5_busy = 1'd0;
reg main_output_8x5_data = 1'd0;
reg [2:0] main_output_8x5_fine_ts = 3'd0;
wire main_output_8x5_override_en;
wire main_output_8x5_override_o;
reg main_output_8x5_previous_data = 1'd0;
wire main_output_8x6_ser_out;
reg [7:0] main_output_8x6_o = 8'd0;
reg main_output_8x6_t_in = 1'd0;
wire main_output_8x6_t_out;
reg main_output_8x6_stb = 1'd0;
reg main_output_8x6_busy = 1'd0;
reg main_output_8x6_data = 1'd0;
reg [2:0] main_output_8x6_fine_ts = 3'd0;
wire main_output_8x6_override_en;
wire main_output_8x6_override_o;
reg main_output_8x6_previous_data = 1'd0;
wire main_output_8x7_ser_out;
reg [7:0] main_output_8x7_o = 8'd0;
reg main_output_8x7_t_in = 1'd0;
wire main_output_8x7_t_out;
reg main_output_8x7_stb = 1'd0;
reg main_output_8x7_busy = 1'd0;
reg main_output_8x7_data = 1'd0;
reg [2:0] main_output_8x7_fine_ts = 3'd0;
wire main_output_8x7_override_en;
wire main_output_8x7_override_o;
reg main_output_8x7_previous_data = 1'd0;
wire main_output_8x8_ser_out;
reg [7:0] main_output_8x8_o = 8'd0;
reg main_output_8x8_t_in = 1'd0;
wire main_output_8x8_t_out;
reg main_output_8x8_stb = 1'd0;
reg main_output_8x8_busy = 1'd0;
reg main_output_8x8_data = 1'd0;
reg [2:0] main_output_8x8_fine_ts = 3'd0;
wire main_output_8x8_override_en;
wire main_output_8x8_override_o;
reg main_output_8x8_previous_data = 1'd0;
wire main_output_8x9_ser_out;
reg [7:0] main_output_8x9_o = 8'd0;
reg main_output_8x9_t_in = 1'd0;
wire main_output_8x9_t_out;
reg main_output_8x9_stb = 1'd0;
reg main_output_8x9_busy = 1'd0;
reg main_output_8x9_data = 1'd0;
reg [2:0] main_output_8x9_fine_ts = 3'd0;
wire main_output_8x9_override_en;
wire main_output_8x9_override_o;
reg main_output_8x9_previous_data = 1'd0;
wire main_output_8x10_ser_out;
reg [7:0] main_output_8x10_o = 8'd0;
reg main_output_8x10_t_in = 1'd0;
wire main_output_8x10_t_out;
reg main_output_8x10_stb = 1'd0;
reg main_output_8x10_busy = 1'd0;
reg main_output_8x10_data = 1'd0;
reg [2:0] main_output_8x10_fine_ts = 3'd0;
wire main_output_8x10_override_en;
wire main_output_8x10_override_o;
reg main_output_8x10_previous_data = 1'd0;
wire main_output_8x11_ser_out;
reg [7:0] main_output_8x11_o = 8'd0;
reg main_output_8x11_t_in = 1'd0;
wire main_output_8x11_t_out;
reg main_output_8x11_stb = 1'd0;
reg main_output_8x11_busy = 1'd0;
reg main_output_8x11_data = 1'd0;
reg [2:0] main_output_8x11_fine_ts = 3'd0;
wire main_output_8x11_override_en;
wire main_output_8x11_override_o;
reg main_output_8x11_previous_data = 1'd0;
wire [2:0] main_spimaster0_interface_cs0;
wire [2:0] main_spimaster0_interface_cs_polarity0;
wire main_spimaster0_interface_clk_next0;
wire main_spimaster0_interface_clk_polarity0;
wire main_spimaster0_interface_cs_next0;
wire main_spimaster0_interface_ce0;
wire main_spimaster0_interface_sample0;
wire main_spimaster0_interface_offline0;
wire main_spimaster0_interface_half_duplex0;
wire main_spimaster0_interface_sdi0;
wire main_spimaster0_interface_sdo0;
reg [2:0] main_spimaster0_interface_cs1 = 3'd7;
reg main_spimaster0_interface_clk0 = 1'd0;
wire main_spimaster0_interface_miso0;
wire main_spimaster0_interface_mosi0;
reg main_spimaster0_interface_miso_reg0 = 1'd0;
reg main_spimaster0_interface_mosi_reg0 = 1'd0;
wire [4:0] main_spimaster0_spimachine0_length0;
wire main_spimaster0_spimachine0_clk_phase0;
reg main_spimaster0_spimachine0_clk_next0;
reg main_spimaster0_spimachine0_cs_next0;
wire main_spimaster0_spimachine0_ce0;
reg main_spimaster0_spimachine0_idle0;
wire main_spimaster0_spimachine0_load0;
reg main_spimaster0_spimachine0_readable0;
reg main_spimaster0_spimachine0_writable0;
wire main_spimaster0_spimachine0_end0;
wire [31:0] main_spimaster0_spimachine0_pdo0;
wire [31:0] main_spimaster0_spimachine0_pdi0;
reg main_spimaster0_spimachine0_sdo0 = 1'd0;
wire main_spimaster0_spimachine0_sdi0;
wire main_spimaster0_spimachine0_lsb_first0;
reg main_spimaster0_spimachine0_load1;
reg main_spimaster0_spimachine0_shift0;
reg main_spimaster0_spimachine0_sample0;
reg [31:0] main_spimaster0_spimachine0_sr0 = 32'd0;
wire [7:0] main_spimaster0_spimachine0_div0;
reg main_spimaster0_spimachine0_extend0;
wire main_spimaster0_spimachine0_done0;
reg main_spimaster0_spimachine0_count0;
reg [6:0] main_spimaster0_spimachine0_cnt0 = 7'd0;
wire main_spimaster0_spimachine0_cnt_done0;
reg main_spimaster0_spimachine0_do_extend0 = 1'd0;
reg [4:0] main_spimaster0_spimachine0_n0 = 5'd0;
reg main_spimaster0_spimachine0_end1 = 1'd0;
reg main_spimaster0_ointerface0_stb0 = 1'd0;
wire main_spimaster0_ointerface0_busy0;
reg [31:0] main_spimaster0_ointerface0_data0 = 32'd0;
reg main_spimaster0_ointerface0_address0 = 1'd0;
wire main_spimaster0_iinterface0_stb0;
wire [31:0] main_spimaster0_iinterface0_data0;
reg main_spimaster0_config_offline0 = 1'd1;
reg main_spimaster0_config_end0 = 1'd1;
reg main_spimaster0_config_input0 = 1'd0;
reg main_spimaster0_config_cs_polarity0 = 1'd0;
reg main_spimaster0_config_clk_polarity0 = 1'd0;
reg main_spimaster0_config_clk_phase0 = 1'd0;
reg main_spimaster0_config_lsb_first0 = 1'd0;
reg main_spimaster0_config_half_duplex0 = 1'd0;
reg [4:0] main_spimaster0_config_length0 = 5'd0;
reg [2:0] main_spimaster0_config_padding0 = 3'd0;
reg [7:0] main_spimaster0_config_div0 = 8'd0;
reg [7:0] main_spimaster0_config_cs0 = 8'd0;
reg main_spimaster0_read0 = 1'd0;
wire main_output_8x0_ser_out1;
reg [7:0] main_output_8x0_o1 = 8'd0;
reg main_output_8x0_t_in1 = 1'd0;
wire main_output_8x0_t_out1;
reg main_output_8x0_stb1 = 1'd0;
reg main_output_8x0_busy1 = 1'd0;
reg main_output_8x0_data1 = 1'd0;
reg [2:0] main_output_8x0_fine_ts1 = 3'd0;
wire main_output_8x0_override_en1;
wire main_output_8x0_override_o1;
reg main_output_8x0_previous_data1 = 1'd0;
reg [31:0] main_urukulmonitor00 = 32'd0;
reg [31:0] main_urukulmonitor01 = 32'd0;
reg [31:0] main_urukulmonitor02 = 32'd0;
reg [31:0] main_urukulmonitor03 = 32'd0;
reg [7:0] main_urukulmonitor0_cs = 8'd0;
reg [31:0] main_urukulmonitor0_current_data = 32'd0;
reg main_urukulmonitor0_current_address = 1'd0;
reg [7:0] main_urukulmonitor0_data_length = 8'd0;
reg [7:0] main_urukulmonitor0_flags = 8'd0;
wire main_urukulmonitor0_ch_sel0;
reg [31:0] main_urukulmonitor0_ftw0 = 32'd0;
wire main_urukulmonitor0_ch_sel1;
reg [31:0] main_urukulmonitor0_ftw1 = 32'd0;
wire main_urukulmonitor0_ch_sel2;
reg [31:0] main_urukulmonitor0_ftw2 = 32'd0;
wire main_urukulmonitor0_ch_sel3;
reg [31:0] main_urukulmonitor0_ftw3 = 32'd0;
wire main_output_8x12_ser_out;
reg [7:0] main_output_8x12_o = 8'd0;
reg main_output_8x12_t_in = 1'd0;
wire main_output_8x12_t_out;
reg main_output_8x12_stb = 1'd0;
reg main_output_8x12_busy = 1'd0;
reg main_output_8x12_data = 1'd0;
reg [2:0] main_output_8x12_fine_ts = 3'd0;
wire main_output_8x12_override_en;
wire main_output_8x12_override_o;
reg main_output_8x12_previous_data = 1'd0;
wire main_output_8x13_ser_out;
reg [7:0] main_output_8x13_o = 8'd0;
reg main_output_8x13_t_in = 1'd0;
wire main_output_8x13_t_out;
reg main_output_8x13_stb = 1'd0;
reg main_output_8x13_busy = 1'd0;
reg main_output_8x13_data = 1'd0;
reg [2:0] main_output_8x13_fine_ts = 3'd0;
wire main_output_8x13_override_en;
wire main_output_8x13_override_o;
reg main_output_8x13_previous_data = 1'd0;
wire main_output_8x14_ser_out;
reg [7:0] main_output_8x14_o = 8'd0;
reg main_output_8x14_t_in = 1'd0;
wire main_output_8x14_t_out;
reg main_output_8x14_stb = 1'd0;
reg main_output_8x14_busy = 1'd0;
reg main_output_8x14_data = 1'd0;
reg [2:0] main_output_8x14_fine_ts = 3'd0;
wire main_output_8x14_override_en;
wire main_output_8x14_override_o;
reg main_output_8x14_previous_data = 1'd0;
wire main_output_8x15_ser_out;
reg [7:0] main_output_8x15_o = 8'd0;
reg main_output_8x15_t_in = 1'd0;
wire main_output_8x15_t_out;
reg main_output_8x15_stb = 1'd0;
reg main_output_8x15_busy = 1'd0;
reg main_output_8x15_data = 1'd0;
reg [2:0] main_output_8x15_fine_ts = 3'd0;
wire main_output_8x15_override_en;
wire main_output_8x15_override_o;
reg main_output_8x15_previous_data = 1'd0;
wire [2:0] main_spimaster1_interface_cs0;
wire [2:0] main_spimaster1_interface_cs_polarity0;
wire main_spimaster1_interface_clk_next0;
wire main_spimaster1_interface_clk_polarity0;
wire main_spimaster1_interface_cs_next0;
wire main_spimaster1_interface_ce0;
wire main_spimaster1_interface_sample0;
wire main_spimaster1_interface_offline0;
wire main_spimaster1_interface_half_duplex0;
wire main_spimaster1_interface_sdi0;
wire main_spimaster1_interface_sdo0;
reg [2:0] main_spimaster1_interface_cs1 = 3'd7;
reg main_spimaster1_interface_clk0 = 1'd0;
wire main_spimaster1_interface_miso0;
wire main_spimaster1_interface_mosi0;
reg main_spimaster1_interface_miso_reg0 = 1'd0;
reg main_spimaster1_interface_mosi_reg0 = 1'd0;
wire [4:0] main_spimaster1_spimachine1_length0;
wire main_spimaster1_spimachine1_clk_phase0;
reg main_spimaster1_spimachine1_clk_next0;
reg main_spimaster1_spimachine1_cs_next0;
wire main_spimaster1_spimachine1_ce0;
reg main_spimaster1_spimachine1_idle0;
wire main_spimaster1_spimachine1_load0;
reg main_spimaster1_spimachine1_readable0;
reg main_spimaster1_spimachine1_writable0;
wire main_spimaster1_spimachine1_end0;
wire [31:0] main_spimaster1_spimachine1_pdo0;
wire [31:0] main_spimaster1_spimachine1_pdi0;
reg main_spimaster1_spimachine1_sdo0 = 1'd0;
wire main_spimaster1_spimachine1_sdi0;
wire main_spimaster1_spimachine1_lsb_first0;
reg main_spimaster1_spimachine1_load1;
reg main_spimaster1_spimachine1_shift0;
reg main_spimaster1_spimachine1_sample0;
reg [31:0] main_spimaster1_spimachine1_sr0 = 32'd0;
wire [7:0] main_spimaster1_spimachine1_div0;
reg main_spimaster1_spimachine1_extend0;
wire main_spimaster1_spimachine1_done0;
reg main_spimaster1_spimachine1_count0;
reg [6:0] main_spimaster1_spimachine1_cnt0 = 7'd0;
wire main_spimaster1_spimachine1_cnt_done0;
reg main_spimaster1_spimachine1_do_extend0 = 1'd0;
reg [4:0] main_spimaster1_spimachine1_n0 = 5'd0;
reg main_spimaster1_spimachine1_end1 = 1'd0;
reg main_spimaster1_ointerface1_stb0 = 1'd0;
wire main_spimaster1_ointerface1_busy0;
reg [31:0] main_spimaster1_ointerface1_data0 = 32'd0;
reg main_spimaster1_ointerface1_address0 = 1'd0;
wire main_spimaster1_iinterface1_stb0;
wire [31:0] main_spimaster1_iinterface1_data0;
reg main_spimaster1_config_offline0 = 1'd1;
reg main_spimaster1_config_end0 = 1'd1;
reg main_spimaster1_config_input0 = 1'd0;
reg main_spimaster1_config_cs_polarity0 = 1'd0;
reg main_spimaster1_config_clk_polarity0 = 1'd0;
reg main_spimaster1_config_clk_phase0 = 1'd0;
reg main_spimaster1_config_lsb_first0 = 1'd0;
reg main_spimaster1_config_half_duplex0 = 1'd0;
reg [4:0] main_spimaster1_config_length0 = 5'd0;
reg [2:0] main_spimaster1_config_padding0 = 3'd0;
reg [7:0] main_spimaster1_config_div0 = 8'd0;
reg [7:0] main_spimaster1_config_cs0 = 8'd0;
reg main_spimaster1_read0 = 1'd0;
wire main_output_8x1_ser_out1;
reg [7:0] main_output_8x1_o1 = 8'd0;
reg main_output_8x1_t_in1 = 1'd0;
wire main_output_8x1_t_out1;
reg main_output_8x1_stb1 = 1'd0;
reg main_output_8x1_busy1 = 1'd0;
reg main_output_8x1_data1 = 1'd0;
reg [2:0] main_output_8x1_fine_ts1 = 3'd0;
wire main_output_8x1_override_en1;
wire main_output_8x1_override_o1;
reg main_output_8x1_previous_data1 = 1'd0;
reg [31:0] main_urukulmonitor10 = 32'd0;
reg [31:0] main_urukulmonitor11 = 32'd0;
reg [31:0] main_urukulmonitor12 = 32'd0;
reg [31:0] main_urukulmonitor13 = 32'd0;
reg [7:0] main_urukulmonitor1_cs = 8'd0;
reg [31:0] main_urukulmonitor1_current_data = 32'd0;
reg main_urukulmonitor1_current_address = 1'd0;
reg [7:0] main_urukulmonitor1_data_length = 8'd0;
reg [7:0] main_urukulmonitor1_flags = 8'd0;
wire main_urukulmonitor1_ch_sel0;
reg [31:0] main_urukulmonitor1_ftw0 = 32'd0;
wire main_urukulmonitor1_ch_sel1;
reg [31:0] main_urukulmonitor1_ftw1 = 32'd0;
wire main_urukulmonitor1_ch_sel2;
reg [31:0] main_urukulmonitor1_ftw2 = 32'd0;
wire main_urukulmonitor1_ch_sel3;
reg [31:0] main_urukulmonitor1_ftw3 = 32'd0;
wire main_output_8x16_ser_out;
reg [7:0] main_output_8x16_o = 8'd0;
reg main_output_8x16_t_in = 1'd0;
wire main_output_8x16_t_out;
reg main_output_8x16_stb = 1'd0;
reg main_output_8x16_busy = 1'd0;
reg main_output_8x16_data = 1'd0;
reg [2:0] main_output_8x16_fine_ts = 3'd0;
wire main_output_8x16_override_en;
wire main_output_8x16_override_o;
reg main_output_8x16_previous_data = 1'd0;
wire main_output_8x17_ser_out;
reg [7:0] main_output_8x17_o = 8'd0;
reg main_output_8x17_t_in = 1'd0;
wire main_output_8x17_t_out;
reg main_output_8x17_stb = 1'd0;
reg main_output_8x17_busy = 1'd0;
reg main_output_8x17_data = 1'd0;
reg [2:0] main_output_8x17_fine_ts = 3'd0;
wire main_output_8x17_override_en;
wire main_output_8x17_override_o;
reg main_output_8x17_previous_data = 1'd0;
wire main_output_8x18_ser_out;
reg [7:0] main_output_8x18_o = 8'd0;
reg main_output_8x18_t_in = 1'd0;
wire main_output_8x18_t_out;
reg main_output_8x18_stb = 1'd0;
reg main_output_8x18_busy = 1'd0;
reg main_output_8x18_data = 1'd0;
reg [2:0] main_output_8x18_fine_ts = 3'd0;
wire main_output_8x18_override_en;
wire main_output_8x18_override_o;
reg main_output_8x18_previous_data = 1'd0;
wire main_output_8x19_ser_out;
reg [7:0] main_output_8x19_o = 8'd0;
reg main_output_8x19_t_in = 1'd0;
wire main_output_8x19_t_out;
reg main_output_8x19_stb = 1'd0;
reg main_output_8x19_busy = 1'd0;
reg main_output_8x19_data = 1'd0;
reg [2:0] main_output_8x19_fine_ts = 3'd0;
wire main_output_8x19_override_en;
wire main_output_8x19_override_o;
reg main_output_8x19_previous_data = 1'd0;
wire main_spimaster0_interface_cs2;
wire main_spimaster0_interface_cs_polarity1;
wire main_spimaster0_interface_clk_next1;
wire main_spimaster0_interface_clk_polarity1;
wire main_spimaster0_interface_cs_next1;
wire main_spimaster0_interface_ce1;
wire main_spimaster0_interface_sample1;
wire main_spimaster0_interface_offline1;
wire main_spimaster0_interface_half_duplex1;
wire main_spimaster0_interface_sdi1;
wire main_spimaster0_interface_sdo1;
reg main_spimaster0_interface_cs3 = 1'd1;
reg main_spimaster0_interface_clk1 = 1'd0;
wire main_spimaster0_interface_miso1;
reg main_spimaster0_interface_mosi1 = 1'd0;
reg main_spimaster0_interface_miso_reg1 = 1'd0;
reg main_spimaster0_interface_mosi_reg1 = 1'd0;
wire [4:0] main_spimaster0_spimachine0_length1;
wire main_spimaster0_spimachine0_clk_phase1;
reg main_spimaster0_spimachine0_clk_next1;
reg main_spimaster0_spimachine0_cs_next1;
wire main_spimaster0_spimachine0_ce1;
reg main_spimaster0_spimachine0_idle1;
wire main_spimaster0_spimachine0_load2;
reg main_spimaster0_spimachine0_readable1;
reg main_spimaster0_spimachine0_writable1;
wire main_spimaster0_spimachine0_end2;
wire [31:0] main_spimaster0_spimachine0_pdo1;
wire [31:0] main_spimaster0_spimachine0_pdi1;
reg main_spimaster0_spimachine0_sdo1 = 1'd0;
wire main_spimaster0_spimachine0_sdi1;
wire main_spimaster0_spimachine0_lsb_first1;
reg main_spimaster0_spimachine0_load3;
reg main_spimaster0_spimachine0_shift1;
reg main_spimaster0_spimachine0_sample1;
reg [31:0] main_spimaster0_spimachine0_sr1 = 32'd0;
wire [7:0] main_spimaster0_spimachine0_div1;
reg main_spimaster0_spimachine0_extend1;
wire main_spimaster0_spimachine0_done1;
reg main_spimaster0_spimachine0_count1;
reg [6:0] main_spimaster0_spimachine0_cnt1 = 7'd0;
wire main_spimaster0_spimachine0_cnt_done1;
reg main_spimaster0_spimachine0_do_extend1 = 1'd0;
reg [4:0] main_spimaster0_spimachine0_n1 = 5'd0;
reg main_spimaster0_spimachine0_end3 = 1'd0;
reg main_spimaster0_ointerface0_stb1 = 1'd0;
wire main_spimaster0_ointerface0_busy1;
reg [31:0] main_spimaster0_ointerface0_data1 = 32'd0;
reg main_spimaster0_ointerface0_address1 = 1'd0;
wire main_spimaster0_iinterface0_stb1;
wire [31:0] main_spimaster0_iinterface0_data1;
reg main_spimaster0_config_offline1 = 1'd1;
reg main_spimaster0_config_end1 = 1'd1;
reg main_spimaster0_config_input1 = 1'd0;
reg main_spimaster0_config_cs_polarity1 = 1'd0;
reg main_spimaster0_config_clk_polarity1 = 1'd0;
reg main_spimaster0_config_clk_phase1 = 1'd0;
reg main_spimaster0_config_lsb_first1 = 1'd0;
reg main_spimaster0_config_half_duplex1 = 1'd0;
reg [4:0] main_spimaster0_config_length1 = 5'd0;
reg [2:0] main_spimaster0_config_padding1 = 3'd0;
reg [7:0] main_spimaster0_config_div1 = 8'd0;
reg [7:0] main_spimaster0_config_cs1 = 8'd0;
reg main_spimaster0_read1 = 1'd0;
wire main_spimaster1_interface_cs2;
wire main_spimaster1_interface_cs_polarity1;
wire main_spimaster1_interface_clk_next1;
wire main_spimaster1_interface_clk_polarity1;
wire main_spimaster1_interface_cs_next1;
wire main_spimaster1_interface_ce1;
wire main_spimaster1_interface_sample1;
wire main_spimaster1_interface_offline1;
wire main_spimaster1_interface_half_duplex1;
wire main_spimaster1_interface_sdi1;
wire main_spimaster1_interface_sdo1;
reg main_spimaster1_interface_cs3 = 1'd1;
reg main_spimaster1_interface_clk1 = 1'd0;
wire main_spimaster1_interface_miso1;
wire main_spimaster1_interface_mosi1;
reg main_spimaster1_interface_miso_reg1 = 1'd0;
reg main_spimaster1_interface_mosi_reg1 = 1'd0;
wire [4:0] main_spimaster1_spimachine1_length1;
wire main_spimaster1_spimachine1_clk_phase1;
reg main_spimaster1_spimachine1_clk_next1;
reg main_spimaster1_spimachine1_cs_next1;
wire main_spimaster1_spimachine1_ce1;
reg main_spimaster1_spimachine1_idle1;
wire main_spimaster1_spimachine1_load2;
reg main_spimaster1_spimachine1_readable1;
reg main_spimaster1_spimachine1_writable1;
wire main_spimaster1_spimachine1_end2;
wire [31:0] main_spimaster1_spimachine1_pdo1;
wire [31:0] main_spimaster1_spimachine1_pdi1;
reg main_spimaster1_spimachine1_sdo1 = 1'd0;
wire main_spimaster1_spimachine1_sdi1;
wire main_spimaster1_spimachine1_lsb_first1;
reg main_spimaster1_spimachine1_load3;
reg main_spimaster1_spimachine1_shift1;
reg main_spimaster1_spimachine1_sample1;
reg [31:0] main_spimaster1_spimachine1_sr1 = 32'd0;
wire [7:0] main_spimaster1_spimachine1_div1;
reg main_spimaster1_spimachine1_extend1;
wire main_spimaster1_spimachine1_done1;
reg main_spimaster1_spimachine1_count1;
reg [6:0] main_spimaster1_spimachine1_cnt1 = 7'd0;
wire main_spimaster1_spimachine1_cnt_done1;
reg main_spimaster1_spimachine1_do_extend1 = 1'd0;
reg [4:0] main_spimaster1_spimachine1_n1 = 5'd0;
reg main_spimaster1_spimachine1_end3 = 1'd0;
reg main_spimaster1_ointerface1_stb1 = 1'd0;
wire main_spimaster1_ointerface1_busy1;
reg [31:0] main_spimaster1_ointerface1_data1 = 32'd0;
reg main_spimaster1_ointerface1_address1 = 1'd0;
wire main_spimaster1_iinterface1_stb1;
wire [31:0] main_spimaster1_iinterface1_data1;
reg main_spimaster1_config_offline1 = 1'd1;
reg main_spimaster1_config_end1 = 1'd1;
reg main_spimaster1_config_input1 = 1'd0;
reg main_spimaster1_config_cs_polarity1 = 1'd0;
reg main_spimaster1_config_clk_polarity1 = 1'd0;
reg main_spimaster1_config_clk_phase1 = 1'd0;
reg main_spimaster1_config_lsb_first1 = 1'd0;
reg main_spimaster1_config_half_duplex1 = 1'd0;
reg [4:0] main_spimaster1_config_length1 = 5'd0;
reg [2:0] main_spimaster1_config_padding1 = 3'd0;
reg [7:0] main_spimaster1_config_div1 = 8'd0;
reg [7:0] main_spimaster1_config_cs1 = 8'd0;
reg main_spimaster1_read1 = 1'd0;
wire main_output_8x20_ser_out;
reg [7:0] main_output_8x20_o = 8'd0;
reg main_output_8x20_t_in = 1'd0;
wire main_output_8x20_t_out;
reg main_output_8x20_stb = 1'd0;
reg main_output_8x20_busy = 1'd0;
reg main_output_8x20_data = 1'd0;
reg [2:0] main_output_8x20_fine_ts = 3'd0;
wire main_output_8x20_override_en;
wire main_output_8x20_override_o;
reg main_output_8x20_previous_data = 1'd0;
wire [1:0] main_spimaster2_interface_cs0;
wire [1:0] main_spimaster2_interface_cs_polarity;
wire main_spimaster2_interface_clk_next;
wire main_spimaster2_interface_clk_polarity;
wire main_spimaster2_interface_cs_next;
wire main_spimaster2_interface_ce;
wire main_spimaster2_interface_sample;
wire main_spimaster2_interface_offline;
wire main_spimaster2_interface_half_duplex;
wire main_spimaster2_interface_sdi;
wire main_spimaster2_interface_sdo;
reg [1:0] main_spimaster2_interface_cs1 = 2'd3;
reg main_spimaster2_interface_clk = 1'd0;
wire main_spimaster2_interface_miso;
wire main_spimaster2_interface_mosi;
reg main_spimaster2_interface_miso_reg = 1'd0;
reg main_spimaster2_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster2_spimachine2_length;
wire main_spimaster2_spimachine2_clk_phase;
reg main_spimaster2_spimachine2_clk_next;
reg main_spimaster2_spimachine2_cs_next;
wire main_spimaster2_spimachine2_ce;
reg main_spimaster2_spimachine2_idle;
wire main_spimaster2_spimachine2_load0;
reg main_spimaster2_spimachine2_readable;
reg main_spimaster2_spimachine2_writable;
wire main_spimaster2_spimachine2_end0;
wire [31:0] main_spimaster2_spimachine2_pdo;
wire [31:0] main_spimaster2_spimachine2_pdi;
reg main_spimaster2_spimachine2_sdo = 1'd0;
wire main_spimaster2_spimachine2_sdi;
wire main_spimaster2_spimachine2_lsb_first;
reg main_spimaster2_spimachine2_load1;
reg main_spimaster2_spimachine2_shift;
reg main_spimaster2_spimachine2_sample;
reg [31:0] main_spimaster2_spimachine2_sr = 32'd0;
wire [7:0] main_spimaster2_spimachine2_div;
reg main_spimaster2_spimachine2_extend;
wire main_spimaster2_spimachine2_done;
reg main_spimaster2_spimachine2_count;
reg [6:0] main_spimaster2_spimachine2_cnt = 7'd0;
wire main_spimaster2_spimachine2_cnt_done;
reg main_spimaster2_spimachine2_do_extend = 1'd0;
reg [4:0] main_spimaster2_spimachine2_n = 5'd0;
reg main_spimaster2_spimachine2_end1 = 1'd0;
reg main_spimaster2_ointerface2_stb = 1'd0;
wire main_spimaster2_ointerface2_busy;
reg [31:0] main_spimaster2_ointerface2_data = 32'd0;
reg main_spimaster2_ointerface2_address = 1'd0;
wire main_spimaster2_iinterface2_stb;
wire [31:0] main_spimaster2_iinterface2_data;
reg main_spimaster2_config_offline = 1'd1;
reg main_spimaster2_config_end = 1'd1;
reg main_spimaster2_config_input = 1'd0;
reg main_spimaster2_config_cs_polarity = 1'd0;
reg main_spimaster2_config_clk_polarity = 1'd0;
reg main_spimaster2_config_clk_phase = 1'd0;
reg main_spimaster2_config_lsb_first = 1'd0;
reg main_spimaster2_config_half_duplex = 1'd0;
reg [4:0] main_spimaster2_config_length = 5'd0;
reg [2:0] main_spimaster2_config_padding = 3'd0;
reg [7:0] main_spimaster2_config_div = 8'd0;
reg [7:0] main_spimaster2_config_cs = 8'd0;
reg main_spimaster2_read = 1'd0;
wire main_ldac_phy_ser_out;
reg [7:0] main_ldac_phy_o = 8'd0;
reg main_ldac_phy_t_in = 1'd0;
wire main_ldac_phy_t_out;
reg main_ldac_phy_stb = 1'd0;
reg main_ldac_phy_busy = 1'd0;
reg main_ldac_phy_data = 1'd0;
reg [2:0] main_ldac_phy_fine_ts = 3'd0;
wire main_ldac_phy_override_en;
wire main_ldac_phy_override_o;
reg main_ldac_phy_previous_data = 1'd0;
wire main_clr_phy_ser_out;
reg [7:0] main_clr_phy_o = 8'd0;
reg main_clr_phy_t_in = 1'd0;
wire main_clr_phy_t_out;
reg main_clr_phy_stb = 1'd0;
reg main_clr_phy_busy = 1'd0;
reg main_clr_phy_data = 1'd0;
reg [2:0] main_clr_phy_fine_ts = 3'd0;
wire main_clr_phy_override_en;
wire main_clr_phy_override_o;
reg main_clr_phy_previous_data = 1'd0;
reg [15:0] main_ad53xxmonitor0 = 16'd0;
reg [15:0] main_ad53xxmonitor1 = 16'd0;
reg [15:0] main_ad53xxmonitor2 = 16'd0;
reg [15:0] main_ad53xxmonitor3 = 16'd0;
reg [15:0] main_ad53xxmonitor4 = 16'd0;
reg [15:0] main_ad53xxmonitor5 = 16'd0;
reg [15:0] main_ad53xxmonitor6 = 16'd0;
reg [15:0] main_ad53xxmonitor7 = 16'd0;
reg [15:0] main_ad53xxmonitor8 = 16'd0;
reg [15:0] main_ad53xxmonitor9 = 16'd0;
reg [15:0] main_ad53xxmonitor10 = 16'd0;
reg [15:0] main_ad53xxmonitor11 = 16'd0;
reg [15:0] main_ad53xxmonitor12 = 16'd0;
reg [15:0] main_ad53xxmonitor13 = 16'd0;
reg [15:0] main_ad53xxmonitor14 = 16'd0;
reg [15:0] main_ad53xxmonitor15 = 16'd0;
reg [15:0] main_ad53xxmonitor16 = 16'd0;
reg [15:0] main_ad53xxmonitor17 = 16'd0;
reg [15:0] main_ad53xxmonitor18 = 16'd0;
reg [15:0] main_ad53xxmonitor19 = 16'd0;
reg [15:0] main_ad53xxmonitor20 = 16'd0;
reg [15:0] main_ad53xxmonitor21 = 16'd0;
reg [15:0] main_ad53xxmonitor22 = 16'd0;
reg [15:0] main_ad53xxmonitor23 = 16'd0;
reg [15:0] main_ad53xxmonitor24 = 16'd0;
reg [15:0] main_ad53xxmonitor25 = 16'd0;
reg [15:0] main_ad53xxmonitor26 = 16'd0;
reg [15:0] main_ad53xxmonitor27 = 16'd0;
reg [15:0] main_ad53xxmonitor28 = 16'd0;
reg [15:0] main_ad53xxmonitor29 = 16'd0;
reg [15:0] main_ad53xxmonitor30 = 16'd0;
reg [15:0] main_ad53xxmonitor31 = 16'd0;
reg [15:0] main_ad53xxmonitor32 = 16'd0;
reg [15:0] main_ad53xxmonitor33 = 16'd0;
reg [15:0] main_ad53xxmonitor34 = 16'd0;
reg [15:0] main_ad53xxmonitor35 = 16'd0;
reg [15:0] main_ad53xxmonitor36 = 16'd0;
reg [15:0] main_ad53xxmonitor37 = 16'd0;
reg [15:0] main_ad53xxmonitor38 = 16'd0;
reg [15:0] main_ad53xxmonitor39 = 16'd0;
reg [15:0] main_ad53xxmonitor40 = 16'd0;
reg [15:0] main_ad53xxmonitor41 = 16'd0;
reg [15:0] main_ad53xxmonitor42 = 16'd0;
reg [15:0] main_ad53xxmonitor43 = 16'd0;
reg [15:0] main_ad53xxmonitor44 = 16'd0;
reg [15:0] main_ad53xxmonitor45 = 16'd0;
reg [15:0] main_ad53xxmonitor46 = 16'd0;
reg [15:0] main_ad53xxmonitor47 = 16'd0;
reg [15:0] main_ad53xxmonitor48 = 16'd0;
reg [15:0] main_ad53xxmonitor49 = 16'd0;
reg [15:0] main_ad53xxmonitor50 = 16'd0;
reg [15:0] main_ad53xxmonitor51 = 16'd0;
reg [15:0] main_ad53xxmonitor52 = 16'd0;
reg [15:0] main_ad53xxmonitor53 = 16'd0;
reg [15:0] main_ad53xxmonitor54 = 16'd0;
reg [15:0] main_ad53xxmonitor55 = 16'd0;
reg [15:0] main_ad53xxmonitor56 = 16'd0;
reg [15:0] main_ad53xxmonitor57 = 16'd0;
reg [15:0] main_ad53xxmonitor58 = 16'd0;
reg [15:0] main_ad53xxmonitor59 = 16'd0;
reg [15:0] main_ad53xxmonitor60 = 16'd0;
reg [15:0] main_ad53xxmonitor61 = 16'd0;
reg [15:0] main_ad53xxmonitor62 = 16'd0;
reg [15:0] main_ad53xxmonitor63 = 16'd0;
reg main_ad53xxmonitor_selected = 1'd0;
reg main_output0_stb = 1'd0;
reg main_output0_busy = 1'd0;
reg main_output0_data = 1'd0;
reg main_output0_pad_o = 1'd0;
wire main_output0_override_en;
wire main_output0_override_o;
reg main_output0_pad_k = 1'd0;
reg main_output1_stb = 1'd0;
reg main_output1_busy = 1'd0;
reg main_output1_data = 1'd0;
reg main_output1_pad_o = 1'd0;
wire main_output1_override_en;
wire main_output1_override_o;
reg main_output1_pad_k = 1'd0;
reg main_output2_stb = 1'd0;
reg main_output2_busy = 1'd0;
reg main_output2_data = 1'd0;
reg main_output2_pad_o = 1'd0;
wire main_output2_override_en;
wire main_output2_override_o;
reg main_output2_pad_k = 1'd0;
reg main_stb = 1'd0;
reg main_busy = 1'd0;
reg [31:0] main_data = 32'd0;
reg [60:0] main_genericstandalone_coarse_ts = 61'd0;
wire [63:0] main_genericstandalone_full_ts;
reg main_genericstandalone_load = 1'd0;
reg [60:0] main_genericstandalone_load_value = 61'd0;
reg [1:0] main_genericstandalone_rtio_core_cri_cmd;
wire [23:0] main_genericstandalone_rtio_core_cri_chan_sel;
wire [63:0] main_genericstandalone_rtio_core_cri_o_timestamp;
wire [511:0] main_genericstandalone_rtio_core_cri_o_data;
wire [7:0] main_genericstandalone_rtio_core_cri_o_address;
wire [2:0] main_genericstandalone_rtio_core_cri_o_status;
reg main_genericstandalone_rtio_core_cri_o_buffer_space_valid = 1'd0;
reg [15:0] main_genericstandalone_rtio_core_cri_o_buffer_space = 16'd0;
wire [63:0] main_genericstandalone_rtio_core_cri_i_timeout;
reg [31:0] main_genericstandalone_rtio_core_cri_i_data = 32'd0;
reg [63:0] main_genericstandalone_rtio_core_cri_i_timestamp = 64'd0;
reg [3:0] main_genericstandalone_rtio_core_cri_i_status = 4'd0;
wire main_genericstandalone_rtio_core_reset_re;
wire main_genericstandalone_rtio_core_reset_r;
reg main_genericstandalone_rtio_core_reset_w = 1'd0;
wire main_genericstandalone_rtio_core_reset_phy_re;
wire main_genericstandalone_rtio_core_reset_phy_r;
reg main_genericstandalone_rtio_core_reset_phy_w = 1'd0;
reg main_genericstandalone_rtio_core_storage_full = 1'd0;
wire main_genericstandalone_rtio_core_storage;
reg main_genericstandalone_rtio_core_re = 1'd0;
wire main_genericstandalone_rtio_core_async_error_re;
wire [2:0] main_genericstandalone_rtio_core_async_error_r;
wire [2:0] main_genericstandalone_rtio_core_async_error_w;
reg [15:0] main_genericstandalone_rtio_core_collision_channel_status = 16'd0;
reg [15:0] main_genericstandalone_rtio_core_busy_channel_status = 16'd0;
reg [15:0] main_genericstandalone_rtio_core_sequence_error_channel_status = 16'd0;
reg main_genericstandalone_rtio_core_cmd_reset = 1'd1;
reg main_genericstandalone_rtio_core_cmd_reset_phy = 1'd1;
wire rio_clk;
wire rio_rst;
wire rio_phy_clk;
wire rio_phy_rst;
reg main_genericstandalone_rtio_core_sed_lane_dist_sequence_error = 1'd0;
reg [15:0] main_genericstandalone_rtio_core_sed_lane_dist_sequence_error_channel = 16'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_minimum_coarse_timestamp = 61'd0;
reg main_genericstandalone_rtio_core_sed_lane_dist_record0_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record0_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record0_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record0_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record1_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record1_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record1_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record1_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record2_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record2_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record2_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record2_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record3_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record3_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record3_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record3_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record4_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record4_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record4_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record4_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record5_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record5_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record5_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record5_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record6_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record6_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record6_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record6_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record7_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record7_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record7_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record7_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record8_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record8_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record8_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record8_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record9_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record9_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record9_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record9_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record10_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record10_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record10_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record10_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record11_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record11_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record11_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record11_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record12_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record12_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record12_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record12_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record13_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record13_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record13_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record13_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record14_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record14_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record14_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record14_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_data;
reg main_genericstandalone_rtio_core_sed_lane_dist_record15_we;
wire main_genericstandalone_rtio_core_sed_lane_dist_record15_writable;
wire main_genericstandalone_rtio_core_sed_lane_dist_record15_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_lane_dist_record15_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_channel;
reg [63:0] main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_data;
wire main_genericstandalone_rtio_core_sed_lane_dist_enable_spread;
wire main_genericstandalone_rtio_core_sed_lane_dist_o_status_wait;
reg main_genericstandalone_rtio_core_sed_lane_dist_o_status_underflow = 1'd0;
reg [3:0] main_genericstandalone_rtio_core_sed_lane_dist_current_lane = 4'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_coarse_timestamp = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps0 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps1 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps2 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps3 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps4 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps5 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps6 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps7 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps8 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps9 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps10 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps11 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps12 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps13 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps14 = 61'd0;
reg [60:0] main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps15 = 61'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_lane_dist_seqn = 13'd0;
wire [60:0] main_genericstandalone_rtio_core_sed_lane_dist_coarse_timestamp;
reg signed [61:0] main_genericstandalone_rtio_core_sed_lane_dist_min_minus_timestamp = 62'sd0;
reg signed [61:0] main_genericstandalone_rtio_core_sed_lane_dist_laneAmin_minus_timestamp = 62'sd0;
reg signed [61:0] main_genericstandalone_rtio_core_sed_lane_dist_laneBmin_minus_timestamp = 62'sd0;
reg signed [61:0] main_genericstandalone_rtio_core_sed_lane_dist_last_minus_timestamp = 62'sd0;
wire [3:0] main_genericstandalone_rtio_core_sed_lane_dist_current_lane_plus_one;
reg main_genericstandalone_rtio_core_sed_lane_dist_quash = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_lane_dist_adr;
wire [13:0] main_genericstandalone_rtio_core_sed_lane_dist_dat_r;
wire signed [13:0] main_genericstandalone_rtio_core_sed_lane_dist_compensation;
wire main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_min;
wire main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_last;
wire main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_laneA_min;
wire main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_laneB_min;
wire main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_lane_min;
reg main_genericstandalone_rtio_core_sed_lane_dist_force_laneB = 1'd0;
reg main_genericstandalone_rtio_core_sed_lane_dist_use_laneB;
reg [3:0] main_genericstandalone_rtio_core_sed_lane_dist_use_lanen;
reg main_genericstandalone_rtio_core_sed_lane_dist_do_write;
reg main_genericstandalone_rtio_core_sed_lane_dist_do_underflow;
reg main_genericstandalone_rtio_core_sed_lane_dist_do_sequence_error;
wire [63:0] main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
wire main_genericstandalone_rtio_core_sed_lane_dist_current_lane_high_watermark;
wire main_genericstandalone_rtio_core_sed_lane_dist_current_lane_writable;
wire main_genericstandalone_rtio_core_sed_record0_we;
wire main_genericstandalone_rtio_core_sed_record0_writable;
wire main_genericstandalone_rtio_core_sed_record0_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record0_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record0_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record0_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record0_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record0_payload_data0;
wire main_genericstandalone_rtio_core_sed_record1_we;
wire main_genericstandalone_rtio_core_sed_record1_writable;
wire main_genericstandalone_rtio_core_sed_record1_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record1_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record1_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record1_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record1_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record1_payload_data0;
wire main_genericstandalone_rtio_core_sed_record2_we;
wire main_genericstandalone_rtio_core_sed_record2_writable;
wire main_genericstandalone_rtio_core_sed_record2_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record2_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record2_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record2_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record2_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record2_payload_data0;
wire main_genericstandalone_rtio_core_sed_record3_we;
wire main_genericstandalone_rtio_core_sed_record3_writable;
wire main_genericstandalone_rtio_core_sed_record3_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record3_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record3_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record3_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record3_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record3_payload_data0;
wire main_genericstandalone_rtio_core_sed_record4_we;
wire main_genericstandalone_rtio_core_sed_record4_writable;
wire main_genericstandalone_rtio_core_sed_record4_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record4_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record4_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record4_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record4_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record4_payload_data0;
wire main_genericstandalone_rtio_core_sed_record5_we;
wire main_genericstandalone_rtio_core_sed_record5_writable;
wire main_genericstandalone_rtio_core_sed_record5_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record5_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record5_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record5_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record5_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record5_payload_data0;
wire main_genericstandalone_rtio_core_sed_record6_we;
wire main_genericstandalone_rtio_core_sed_record6_writable;
wire main_genericstandalone_rtio_core_sed_record6_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record6_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record6_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record6_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record6_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record6_payload_data0;
wire main_genericstandalone_rtio_core_sed_record7_we;
wire main_genericstandalone_rtio_core_sed_record7_writable;
wire main_genericstandalone_rtio_core_sed_record7_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record7_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record7_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record7_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record7_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record7_payload_data0;
wire main_genericstandalone_rtio_core_sed_record8_we;
wire main_genericstandalone_rtio_core_sed_record8_writable;
wire main_genericstandalone_rtio_core_sed_record8_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record8_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record8_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record8_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record8_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record8_payload_data0;
wire main_genericstandalone_rtio_core_sed_record9_we;
wire main_genericstandalone_rtio_core_sed_record9_writable;
wire main_genericstandalone_rtio_core_sed_record9_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record9_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record9_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record9_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record9_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record9_payload_data0;
wire main_genericstandalone_rtio_core_sed_record10_we;
wire main_genericstandalone_rtio_core_sed_record10_writable;
wire main_genericstandalone_rtio_core_sed_record10_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record10_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record10_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record10_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record10_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record10_payload_data0;
wire main_genericstandalone_rtio_core_sed_record11_we;
wire main_genericstandalone_rtio_core_sed_record11_writable;
wire main_genericstandalone_rtio_core_sed_record11_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record11_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record11_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record11_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record11_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record11_payload_data0;
wire main_genericstandalone_rtio_core_sed_record12_we;
wire main_genericstandalone_rtio_core_sed_record12_writable;
wire main_genericstandalone_rtio_core_sed_record12_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record12_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record12_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record12_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record12_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record12_payload_data0;
wire main_genericstandalone_rtio_core_sed_record13_we;
wire main_genericstandalone_rtio_core_sed_record13_writable;
wire main_genericstandalone_rtio_core_sed_record13_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record13_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record13_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record13_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record13_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record13_payload_data0;
wire main_genericstandalone_rtio_core_sed_record14_we;
wire main_genericstandalone_rtio_core_sed_record14_writable;
wire main_genericstandalone_rtio_core_sed_record14_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record14_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record14_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record14_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record14_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record14_payload_data0;
wire main_genericstandalone_rtio_core_sed_record15_we;
wire main_genericstandalone_rtio_core_sed_record15_writable;
wire main_genericstandalone_rtio_core_sed_record15_high_watermark;
wire [12:0] main_genericstandalone_rtio_core_sed_record15_seqn0;
wire [5:0] main_genericstandalone_rtio_core_sed_record15_payload_channel0;
wire [63:0] main_genericstandalone_rtio_core_sed_record15_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record15_payload_address0;
wire [31:0] main_genericstandalone_rtio_core_sed_record15_payload_data0;
wire main_genericstandalone_rtio_core_sed_record16_re;
wire main_genericstandalone_rtio_core_sed_record16_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record16_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record16_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record16_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record16_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record16_payload_data;
wire main_genericstandalone_rtio_core_sed_record17_re;
wire main_genericstandalone_rtio_core_sed_record17_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record17_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record17_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record17_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record17_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record17_payload_data;
wire main_genericstandalone_rtio_core_sed_record18_re;
wire main_genericstandalone_rtio_core_sed_record18_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record18_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record18_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record18_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record18_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record18_payload_data;
wire main_genericstandalone_rtio_core_sed_record19_re;
wire main_genericstandalone_rtio_core_sed_record19_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record19_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record19_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record19_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record19_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record19_payload_data;
wire main_genericstandalone_rtio_core_sed_record20_re;
wire main_genericstandalone_rtio_core_sed_record20_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record20_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record20_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record20_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record20_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record20_payload_data;
wire main_genericstandalone_rtio_core_sed_record21_re;
wire main_genericstandalone_rtio_core_sed_record21_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record21_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record21_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record21_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record21_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record21_payload_data;
wire main_genericstandalone_rtio_core_sed_record22_re;
wire main_genericstandalone_rtio_core_sed_record22_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record22_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record22_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record22_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record22_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record22_payload_data;
wire main_genericstandalone_rtio_core_sed_record23_re;
wire main_genericstandalone_rtio_core_sed_record23_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record23_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record23_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record23_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record23_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record23_payload_data;
wire main_genericstandalone_rtio_core_sed_record24_re;
wire main_genericstandalone_rtio_core_sed_record24_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record24_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record24_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record24_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record24_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record24_payload_data;
wire main_genericstandalone_rtio_core_sed_record25_re;
wire main_genericstandalone_rtio_core_sed_record25_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record25_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record25_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record25_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record25_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record25_payload_data;
wire main_genericstandalone_rtio_core_sed_record26_re;
wire main_genericstandalone_rtio_core_sed_record26_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record26_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record26_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record26_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record26_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record26_payload_data;
wire main_genericstandalone_rtio_core_sed_record27_re;
wire main_genericstandalone_rtio_core_sed_record27_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record27_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record27_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record27_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record27_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record27_payload_data;
wire main_genericstandalone_rtio_core_sed_record28_re;
wire main_genericstandalone_rtio_core_sed_record28_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record28_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record28_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record28_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record28_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record28_payload_data;
wire main_genericstandalone_rtio_core_sed_record29_re;
wire main_genericstandalone_rtio_core_sed_record29_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record29_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record29_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record29_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record29_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record29_payload_data;
wire main_genericstandalone_rtio_core_sed_record30_re;
wire main_genericstandalone_rtio_core_sed_record30_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record30_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record30_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record30_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record30_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record30_payload_data;
wire main_genericstandalone_rtio_core_sed_record31_re;
wire main_genericstandalone_rtio_core_sed_record31_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_record31_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_record31_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_record31_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_record31_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_record31_payload_data;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered0_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered0_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered0_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered0_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered0_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered1_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered1_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered1_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered1_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered1_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered2_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered2_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered2_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered2_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered2_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered3_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered3_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered3_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered3_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered3_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered4_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered4_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered4_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered4_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered4_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered5_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered5_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered5_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered5_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered5_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered6_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered6_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered6_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered6_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered6_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered7_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered7_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered7_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered7_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered7_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered8_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered8_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered8_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered8_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered8_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered9_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered9_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered9_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered9_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered9_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered10_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered10_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered10_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered10_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered10_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered11_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered11_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered11_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered11_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered11_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered12_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered12_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered12_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered12_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered12_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered13_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered13_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered13_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered13_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered13_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered14_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered14_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered14_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered14_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered14_level1;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered15_re;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered15_readable = 1'd0;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_we;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_writable;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_re;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_readable;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_din;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_dout;
reg [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 = 8'd0;
reg main_genericstandalone_rtio_core_sed_syncfifobuffered15_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_we;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_dat_w;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered15_do_read;
wire [6:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_adr;
wire [116:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_dat_r;
wire main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_re;
wire [7:0] main_genericstandalone_rtio_core_sed_syncfifobuffered15_level1;
wire main_genericstandalone_rtio_core_sed_gates_record0_re;
wire main_genericstandalone_rtio_core_sed_gates_record0_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record0_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record0_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record0_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record0_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record0_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record1_re;
wire main_genericstandalone_rtio_core_sed_gates_record1_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record1_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record1_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record1_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record1_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record1_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record2_re;
wire main_genericstandalone_rtio_core_sed_gates_record2_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record2_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record2_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record2_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record2_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record2_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record3_re;
wire main_genericstandalone_rtio_core_sed_gates_record3_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record3_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record3_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record3_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record3_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record3_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record4_re;
wire main_genericstandalone_rtio_core_sed_gates_record4_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record4_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record4_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record4_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record4_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record4_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record5_re;
wire main_genericstandalone_rtio_core_sed_gates_record5_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record5_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record5_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record5_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record5_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record5_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record6_re;
wire main_genericstandalone_rtio_core_sed_gates_record6_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record6_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record6_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record6_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record6_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record6_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record7_re;
wire main_genericstandalone_rtio_core_sed_gates_record7_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record7_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record7_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record7_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record7_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record7_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record8_re;
wire main_genericstandalone_rtio_core_sed_gates_record8_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record8_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record8_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record8_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record8_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record8_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record9_re;
wire main_genericstandalone_rtio_core_sed_gates_record9_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record9_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record9_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record9_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record9_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record9_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record10_re;
wire main_genericstandalone_rtio_core_sed_gates_record10_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record10_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record10_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record10_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record10_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record10_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record11_re;
wire main_genericstandalone_rtio_core_sed_gates_record11_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record11_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record11_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record11_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record11_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record11_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record12_re;
wire main_genericstandalone_rtio_core_sed_gates_record12_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record12_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record12_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record12_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record12_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record12_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record13_re;
wire main_genericstandalone_rtio_core_sed_gates_record13_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record13_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record13_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record13_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record13_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record13_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record14_re;
wire main_genericstandalone_rtio_core_sed_gates_record14_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record14_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record14_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record14_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record14_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record14_payload_data;
wire main_genericstandalone_rtio_core_sed_gates_record15_re;
wire main_genericstandalone_rtio_core_sed_gates_record15_readable;
wire [12:0] main_genericstandalone_rtio_core_sed_gates_record15_seqn;
wire [5:0] main_genericstandalone_rtio_core_sed_gates_record15_payload_channel;
wire [63:0] main_genericstandalone_rtio_core_sed_gates_record15_payload_timestamp;
wire [1:0] main_genericstandalone_rtio_core_sed_gates_record15_payload_address;
wire [31:0] main_genericstandalone_rtio_core_sed_gates_record15_payload_data;
reg main_genericstandalone_rtio_core_sed_gates_record16_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record16_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record16_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record16_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record16_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record16_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record16_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record16_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record17_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record17_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record17_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record17_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record17_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record17_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record17_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record17_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record18_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record18_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record18_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record18_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record18_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record18_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record18_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record18_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record19_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record19_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record19_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record19_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record19_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record19_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record19_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record19_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record20_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record20_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record20_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record20_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record20_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record20_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record20_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record20_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record21_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record21_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record21_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record21_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record21_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record21_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record21_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record21_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record22_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record22_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record22_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record22_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record22_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record22_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record22_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record22_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record23_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record23_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record23_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record23_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record23_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record23_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record23_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record23_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record24_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record24_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record24_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record24_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record24_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record24_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record24_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record24_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record25_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record25_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record25_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record25_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record25_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record25_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record25_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record25_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record26_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record26_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record26_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record26_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record26_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record26_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record26_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record26_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record27_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record27_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record27_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record27_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record27_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record27_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record27_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record27_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record28_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record28_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record28_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record28_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record28_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record28_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record28_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record28_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record29_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record29_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record29_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record29_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record29_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record29_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record29_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record29_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record30_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record30_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record30_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record30_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record30_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record30_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record30_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record30_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_gates_record31_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_gates_record31_seqn = 13'd0;
wire main_genericstandalone_rtio_core_sed_gates_record31_replace_occured;
wire main_genericstandalone_rtio_core_sed_gates_record31_nondata_replace_occured;
reg [5:0] main_genericstandalone_rtio_core_sed_gates_record31_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_gates_record31_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_gates_record31_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_gates_record31_payload_data = 32'd0;
wire [60:0] main_genericstandalone_rtio_core_sed_gates_coarse_timestamp;
reg main_genericstandalone_rtio_core_sed_collision = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_collision_channel = 6'd0;
reg main_genericstandalone_rtio_core_sed_busy = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_busy_channel = 6'd0;
wire main_genericstandalone_rtio_core_sed_record0_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record0_seqn1;
wire main_genericstandalone_rtio_core_sed_record0_replace_occured;
wire main_genericstandalone_rtio_core_sed_record0_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record0_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record0_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record0_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record0_payload_data1;
wire main_genericstandalone_rtio_core_sed_record1_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record1_seqn1;
wire main_genericstandalone_rtio_core_sed_record1_replace_occured;
wire main_genericstandalone_rtio_core_sed_record1_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record1_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record1_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record1_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record1_payload_data1;
wire main_genericstandalone_rtio_core_sed_record2_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record2_seqn1;
wire main_genericstandalone_rtio_core_sed_record2_replace_occured;
wire main_genericstandalone_rtio_core_sed_record2_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record2_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record2_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record2_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record2_payload_data1;
wire main_genericstandalone_rtio_core_sed_record3_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record3_seqn1;
wire main_genericstandalone_rtio_core_sed_record3_replace_occured;
wire main_genericstandalone_rtio_core_sed_record3_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record3_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record3_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record3_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record3_payload_data1;
wire main_genericstandalone_rtio_core_sed_record4_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record4_seqn1;
wire main_genericstandalone_rtio_core_sed_record4_replace_occured;
wire main_genericstandalone_rtio_core_sed_record4_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record4_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record4_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record4_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record4_payload_data1;
wire main_genericstandalone_rtio_core_sed_record5_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record5_seqn1;
wire main_genericstandalone_rtio_core_sed_record5_replace_occured;
wire main_genericstandalone_rtio_core_sed_record5_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record5_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record5_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record5_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record5_payload_data1;
wire main_genericstandalone_rtio_core_sed_record6_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record6_seqn1;
wire main_genericstandalone_rtio_core_sed_record6_replace_occured;
wire main_genericstandalone_rtio_core_sed_record6_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record6_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record6_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record6_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record6_payload_data1;
wire main_genericstandalone_rtio_core_sed_record7_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record7_seqn1;
wire main_genericstandalone_rtio_core_sed_record7_replace_occured;
wire main_genericstandalone_rtio_core_sed_record7_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record7_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record7_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record7_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record7_payload_data1;
wire main_genericstandalone_rtio_core_sed_record8_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record8_seqn1;
wire main_genericstandalone_rtio_core_sed_record8_replace_occured;
wire main_genericstandalone_rtio_core_sed_record8_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record8_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record8_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record8_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record8_payload_data1;
wire main_genericstandalone_rtio_core_sed_record9_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record9_seqn1;
wire main_genericstandalone_rtio_core_sed_record9_replace_occured;
wire main_genericstandalone_rtio_core_sed_record9_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record9_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record9_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record9_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record9_payload_data1;
wire main_genericstandalone_rtio_core_sed_record10_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record10_seqn1;
wire main_genericstandalone_rtio_core_sed_record10_replace_occured;
wire main_genericstandalone_rtio_core_sed_record10_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record10_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record10_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record10_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record10_payload_data1;
wire main_genericstandalone_rtio_core_sed_record11_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record11_seqn1;
wire main_genericstandalone_rtio_core_sed_record11_replace_occured;
wire main_genericstandalone_rtio_core_sed_record11_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record11_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record11_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record11_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record11_payload_data1;
wire main_genericstandalone_rtio_core_sed_record12_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record12_seqn1;
wire main_genericstandalone_rtio_core_sed_record12_replace_occured;
wire main_genericstandalone_rtio_core_sed_record12_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record12_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record12_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record12_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record12_payload_data1;
wire main_genericstandalone_rtio_core_sed_record13_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record13_seqn1;
wire main_genericstandalone_rtio_core_sed_record13_replace_occured;
wire main_genericstandalone_rtio_core_sed_record13_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record13_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record13_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record13_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record13_payload_data1;
wire main_genericstandalone_rtio_core_sed_record14_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record14_seqn1;
wire main_genericstandalone_rtio_core_sed_record14_replace_occured;
wire main_genericstandalone_rtio_core_sed_record14_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record14_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record14_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record14_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record14_payload_data1;
wire main_genericstandalone_rtio_core_sed_record15_valid0;
wire [12:0] main_genericstandalone_rtio_core_sed_record15_seqn1;
wire main_genericstandalone_rtio_core_sed_record15_replace_occured;
wire main_genericstandalone_rtio_core_sed_record15_nondata_replace_occured;
wire [5:0] main_genericstandalone_rtio_core_sed_record15_payload_channel1;
wire [2:0] main_genericstandalone_rtio_core_sed_record15_payload_fine_ts0;
wire [1:0] main_genericstandalone_rtio_core_sed_record15_payload_address1;
wire [31:0] main_genericstandalone_rtio_core_sed_record15_payload_data1;
reg main_genericstandalone_rtio_core_sed_record0_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record0_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record0_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record0_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record0_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record0_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record1_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record1_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record1_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record1_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record1_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record1_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record2_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record2_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record2_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record2_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record2_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record2_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record3_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record3_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record3_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record3_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record3_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record3_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record4_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record4_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record4_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record4_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record4_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record4_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record5_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record5_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record5_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record5_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record5_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record5_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record6_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record6_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record6_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record6_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record6_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record6_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record7_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record7_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record7_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record7_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record7_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record7_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record8_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record8_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record8_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record8_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record8_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record8_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record9_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record9_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record9_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record9_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record9_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record9_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record10_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record10_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record10_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record10_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record10_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record10_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record11_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record11_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record11_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record11_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record11_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record11_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record12_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record12_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record12_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record12_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record12_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record12_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record13_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record13_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record13_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record13_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record13_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record13_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record14_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record14_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record14_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record14_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record14_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record14_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record15_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record15_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record15_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record15_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record15_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record15_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference0;
reg main_genericstandalone_rtio_core_sed_nondata_difference1;
reg main_genericstandalone_rtio_core_sed_nondata_difference2;
reg main_genericstandalone_rtio_core_sed_nondata_difference3;
reg main_genericstandalone_rtio_core_sed_nondata_difference4;
reg main_genericstandalone_rtio_core_sed_nondata_difference5;
reg main_genericstandalone_rtio_core_sed_nondata_difference6;
reg main_genericstandalone_rtio_core_sed_nondata_difference7;
reg main_genericstandalone_rtio_core_sed_record16_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record16_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record16_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record16_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record16_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record16_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record16_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record16_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record17_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record17_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record17_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record17_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record17_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record17_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record18_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record18_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record18_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record18_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record18_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record18_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record19_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record19_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record19_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record19_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record19_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record19_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record19_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record19_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record20_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record20_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record20_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record20_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record20_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record20_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record20_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record20_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record21_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record21_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record21_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record21_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record21_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record21_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record22_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record22_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record22_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record22_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record22_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record22_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record23_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record23_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record23_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record23_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record23_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record23_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record23_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record23_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record24_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record24_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record24_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record24_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record24_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record24_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record24_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record24_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record25_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record25_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record25_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record25_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record25_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record25_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record26_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record26_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record26_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record26_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record26_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record26_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record27_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record27_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record27_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record27_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record27_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record27_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record27_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record27_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record28_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record28_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record28_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record28_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record28_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record28_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record28_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record28_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record29_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record29_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record29_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record29_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record29_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record29_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record30_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record30_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record30_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record30_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record30_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record30_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record31_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record31_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record31_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record31_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record31_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record31_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record31_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record31_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference8;
reg main_genericstandalone_rtio_core_sed_nondata_difference9;
reg main_genericstandalone_rtio_core_sed_nondata_difference10;
reg main_genericstandalone_rtio_core_sed_nondata_difference11;
reg main_genericstandalone_rtio_core_sed_nondata_difference12;
reg main_genericstandalone_rtio_core_sed_nondata_difference13;
reg main_genericstandalone_rtio_core_sed_nondata_difference14;
reg main_genericstandalone_rtio_core_sed_nondata_difference15;
reg main_genericstandalone_rtio_core_sed_record32_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record32_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record32_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record32_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record32_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record32_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record32_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record32_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record33_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record33_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record33_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record33_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record33_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record33_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record34_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record34_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record34_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record34_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record34_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record34_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record35_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record35_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record35_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record35_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record35_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record35_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record35_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record35_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record36_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record36_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record36_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record36_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record36_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record36_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record36_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record36_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record37_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record37_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record37_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record37_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record37_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record37_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record38_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record38_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record38_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record38_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record38_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record38_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record39_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record39_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record39_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record39_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record39_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record39_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record39_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record39_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record40_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record40_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record40_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record40_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record40_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record40_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record40_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record40_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record41_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record41_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record41_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record41_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record41_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record41_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record42_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record42_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record42_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record42_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record42_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record42_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record43_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record43_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record43_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record43_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record43_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record43_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record43_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record43_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record44_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record44_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record44_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record44_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record44_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record44_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record44_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record44_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record45_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record45_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record45_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record45_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record45_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record45_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record46_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record46_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record46_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record46_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record46_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record46_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record47_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record47_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record47_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record47_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record47_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record47_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record47_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record47_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference16;
reg main_genericstandalone_rtio_core_sed_nondata_difference17;
reg main_genericstandalone_rtio_core_sed_nondata_difference18;
reg main_genericstandalone_rtio_core_sed_nondata_difference19;
reg main_genericstandalone_rtio_core_sed_record48_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record48_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record48_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record48_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record48_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record48_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record48_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record48_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record49_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record49_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record49_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record49_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record49_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record49_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record49_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record49_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record50_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record50_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record50_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record50_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record50_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record50_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record51_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record51_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record51_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record51_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record51_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record51_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record52_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record52_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record52_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record52_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record52_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record52_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record53_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record53_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record53_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record53_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record53_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record53_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record54_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record54_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record54_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record54_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record54_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record54_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record54_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record54_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record55_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record55_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record55_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record55_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record55_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record55_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record55_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record55_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record56_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record56_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record56_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record56_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record56_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record56_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record56_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record56_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record57_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record57_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record57_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record57_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record57_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record57_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record57_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record57_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record58_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record58_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record58_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record58_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record58_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record58_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record59_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record59_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record59_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record59_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record59_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record59_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record60_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record60_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record60_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record60_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record60_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record60_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record61_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record61_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record61_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record61_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record61_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record61_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record62_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record62_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record62_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record62_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record62_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record62_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record62_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record62_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record63_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record63_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record63_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record63_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record63_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record63_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record63_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record63_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference20;
reg main_genericstandalone_rtio_core_sed_nondata_difference21;
reg main_genericstandalone_rtio_core_sed_nondata_difference22;
reg main_genericstandalone_rtio_core_sed_nondata_difference23;
reg main_genericstandalone_rtio_core_sed_nondata_difference24;
reg main_genericstandalone_rtio_core_sed_nondata_difference25;
reg main_genericstandalone_rtio_core_sed_nondata_difference26;
reg main_genericstandalone_rtio_core_sed_nondata_difference27;
reg main_genericstandalone_rtio_core_sed_record64_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record64_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record64_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record64_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record64_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record64_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record64_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record64_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record65_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record65_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record65_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record65_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record65_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record65_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record65_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record65_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record66_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record66_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record66_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record66_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record66_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record66_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record67_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record67_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record67_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record67_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record67_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record67_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record68_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record68_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record68_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record68_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record68_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record68_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record69_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record69_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record69_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record69_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record69_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record69_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record70_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record70_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record70_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record70_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record70_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record70_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record70_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record70_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record71_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record71_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record71_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record71_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record71_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record71_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record71_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record71_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record72_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record72_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record72_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record72_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record72_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record72_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record72_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record72_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record73_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record73_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record73_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record73_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record73_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record73_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record73_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record73_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record74_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record74_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record74_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record74_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record74_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record74_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record75_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record75_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record75_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record75_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record75_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record75_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record76_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record76_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record76_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record76_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record76_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record76_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record77_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record77_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record77_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record77_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record77_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record77_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record78_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record78_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record78_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record78_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record78_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record78_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record78_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record78_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record79_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record79_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record79_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record79_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record79_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record79_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record79_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record79_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference28;
reg main_genericstandalone_rtio_core_sed_nondata_difference29;
reg main_genericstandalone_rtio_core_sed_nondata_difference30;
reg main_genericstandalone_rtio_core_sed_nondata_difference31;
reg main_genericstandalone_rtio_core_sed_record80_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record80_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record80_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record80_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record80_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record80_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record80_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record80_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record81_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record81_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record81_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record81_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record81_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record81_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record82_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record82_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record82_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record82_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record82_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record82_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record83_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record83_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record83_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record83_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record83_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record83_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record84_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record84_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record84_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record84_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record84_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record84_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record85_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record85_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record85_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record85_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record85_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record85_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record86_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record86_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record86_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record86_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record86_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record86_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record87_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record87_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record87_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record87_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record87_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record87_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record87_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record87_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record88_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record88_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record88_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record88_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record88_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record88_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record88_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record88_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record89_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record89_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record89_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record89_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record89_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record89_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record90_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record90_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record90_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record90_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record90_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record90_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record91_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record91_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record91_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record91_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record91_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record91_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record92_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record92_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record92_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record92_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record92_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record92_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record93_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record93_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record93_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record93_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record93_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record93_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record94_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record94_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record94_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record94_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record94_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record94_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record95_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record95_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record95_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record95_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record95_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record95_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record95_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record95_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference32;
reg main_genericstandalone_rtio_core_sed_nondata_difference33;
reg main_genericstandalone_rtio_core_sed_nondata_difference34;
reg main_genericstandalone_rtio_core_sed_nondata_difference35;
reg main_genericstandalone_rtio_core_sed_nondata_difference36;
reg main_genericstandalone_rtio_core_sed_nondata_difference37;
reg main_genericstandalone_rtio_core_sed_record96_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record96_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record96_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record96_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record96_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record96_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record96_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record96_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record97_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record97_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record97_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record97_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record97_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record97_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record97_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record97_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record98_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record98_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record98_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record98_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record98_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record98_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record98_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record98_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record99_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record99_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record99_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record99_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record99_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record99_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record99_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record99_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record100_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record100_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record100_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record100_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record100_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record100_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record101_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record101_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record101_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record101_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record101_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record101_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record102_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record102_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record102_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record102_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record102_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record102_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record103_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record103_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record103_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record103_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record103_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record103_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record104_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record104_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record104_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record104_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record104_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record104_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record105_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record105_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record105_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record105_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record105_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record105_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record106_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record106_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record106_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record106_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record106_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record106_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record107_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record107_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record107_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record107_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record107_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record107_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record108_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record108_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record108_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record108_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record108_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record108_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record108_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record108_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record109_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record109_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record109_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record109_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record109_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record109_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record109_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record109_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record110_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record110_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record110_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record110_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record110_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record110_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record110_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record110_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record111_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record111_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record111_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record111_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record111_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record111_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record111_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record111_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference38;
reg main_genericstandalone_rtio_core_sed_nondata_difference39;
reg main_genericstandalone_rtio_core_sed_nondata_difference40;
reg main_genericstandalone_rtio_core_sed_nondata_difference41;
reg main_genericstandalone_rtio_core_sed_nondata_difference42;
reg main_genericstandalone_rtio_core_sed_nondata_difference43;
reg main_genericstandalone_rtio_core_sed_nondata_difference44;
reg main_genericstandalone_rtio_core_sed_nondata_difference45;
reg main_genericstandalone_rtio_core_sed_record112_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record112_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record112_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record112_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record112_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record112_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record112_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record112_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record113_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record113_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record113_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record113_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record113_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record113_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record113_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record113_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record114_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record114_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record114_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record114_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record114_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record114_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record114_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record114_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record115_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record115_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record115_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record115_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record115_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record115_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record115_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record115_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record116_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record116_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record116_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record116_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record116_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record116_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record117_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record117_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record117_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record117_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record117_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record117_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record118_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record118_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record118_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record118_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record118_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record118_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record119_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record119_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record119_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record119_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record119_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record119_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record120_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record120_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record120_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record120_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record120_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record120_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record121_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record121_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record121_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record121_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record121_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record121_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record122_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record122_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record122_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record122_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record122_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record122_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record123_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record123_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record123_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record123_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record123_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record123_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record124_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record124_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record124_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record124_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record124_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record124_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record124_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record124_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record125_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record125_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record125_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record125_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record125_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record125_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record125_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record125_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record126_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record126_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record126_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record126_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record126_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record126_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record126_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record126_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record127_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record127_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record127_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record127_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record127_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record127_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record127_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record127_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference46;
reg main_genericstandalone_rtio_core_sed_nondata_difference47;
reg main_genericstandalone_rtio_core_sed_nondata_difference48;
reg main_genericstandalone_rtio_core_sed_nondata_difference49;
reg main_genericstandalone_rtio_core_sed_record128_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record128_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record128_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record128_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record128_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record128_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record128_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record128_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record129_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record129_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record129_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record129_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record129_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record129_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record129_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record129_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record130_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record130_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record130_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record130_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record130_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record130_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record131_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record131_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record131_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record131_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record131_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record131_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record132_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record132_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record132_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record132_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record132_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record132_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record133_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record133_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record133_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record133_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record133_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record133_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record134_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record134_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record134_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record134_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record134_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record134_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record135_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record135_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record135_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record135_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record135_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record135_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record136_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record136_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record136_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record136_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record136_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record136_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record137_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record137_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record137_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record137_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record137_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record137_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record138_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record138_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record138_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record138_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record138_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record138_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record139_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record139_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record139_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record139_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record139_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record139_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record140_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record140_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record140_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record140_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record140_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record140_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record141_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record141_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record141_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record141_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record141_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record141_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record142_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record142_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record142_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record142_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record142_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record142_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record142_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record142_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record143_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record143_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record143_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record143_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record143_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record143_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record143_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record143_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference50;
reg main_genericstandalone_rtio_core_sed_nondata_difference51;
reg main_genericstandalone_rtio_core_sed_nondata_difference52;
reg main_genericstandalone_rtio_core_sed_nondata_difference53;
reg main_genericstandalone_rtio_core_sed_nondata_difference54;
reg main_genericstandalone_rtio_core_sed_nondata_difference55;
reg main_genericstandalone_rtio_core_sed_record144_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record144_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record144_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record144_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record144_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record144_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record144_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record144_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record145_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record145_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record145_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record145_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record145_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record145_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record145_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record145_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record146_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record146_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record146_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record146_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record146_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record146_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record146_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record146_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record147_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record147_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record147_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record147_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record147_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record147_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record147_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record147_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record148_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record148_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record148_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record148_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record148_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record148_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record148_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record148_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record149_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record149_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record149_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record149_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record149_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record149_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record149_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record149_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record150_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record150_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record150_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record150_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record150_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record150_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record150_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record150_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record151_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record151_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record151_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record151_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record151_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record151_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record151_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record151_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record152_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record152_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record152_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record152_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record152_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record152_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record152_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record152_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record153_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record153_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record153_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record153_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record153_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record153_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record153_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record153_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record154_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record154_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record154_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record154_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record154_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record154_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record154_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record154_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record155_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record155_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record155_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record155_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record155_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record155_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record155_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record155_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record156_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record156_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record156_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record156_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record156_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record156_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record156_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record156_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record157_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record157_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record157_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record157_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record157_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record157_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record157_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record157_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record158_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record158_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record158_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record158_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record158_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record158_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record158_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record158_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_record159_rec_valid = 1'd0;
reg [12:0] main_genericstandalone_rtio_core_sed_record159_rec_seqn = 13'd0;
reg main_genericstandalone_rtio_core_sed_record159_rec_replace_occured = 1'd0;
reg main_genericstandalone_rtio_core_sed_record159_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_record159_rec_payload_channel = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record159_rec_payload_fine_ts = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record159_rec_payload_address = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record159_rec_payload_data = 32'd0;
reg main_genericstandalone_rtio_core_sed_nondata_difference56;
reg main_genericstandalone_rtio_core_sed_nondata_difference57;
reg main_genericstandalone_rtio_core_sed_nondata_difference58;
reg main_genericstandalone_rtio_core_sed_nondata_difference59;
reg main_genericstandalone_rtio_core_sed_nondata_difference60;
reg main_genericstandalone_rtio_core_sed_nondata_difference61;
reg main_genericstandalone_rtio_core_sed_nondata_difference62;
reg main_genericstandalone_rtio_core_sed_record0_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record0_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record0_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record0_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record0_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record1_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record1_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record1_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record1_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record1_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record2_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record2_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record2_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record2_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record2_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record3_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record3_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record3_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record3_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record3_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record4_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record4_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record4_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record4_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record4_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record5_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record5_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record5_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record5_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record5_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record6_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record6_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record6_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record6_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record6_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record7_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record7_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record7_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record7_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record7_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record8_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record8_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record8_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record8_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record8_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record9_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record9_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record9_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record9_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record9_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record10_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record10_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record10_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record10_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record10_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record11_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record11_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record11_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record11_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record11_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record12_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record12_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record12_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record12_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record12_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record13_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record13_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record13_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record13_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record13_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record14_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record14_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record14_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record14_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record14_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_record15_valid1 = 1'd0;
wire main_genericstandalone_rtio_core_sed_record15_collision;
reg [5:0] main_genericstandalone_rtio_core_sed_record15_payload_channel2 = 6'd0;
reg [2:0] main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1 = 3'd0;
reg [1:0] main_genericstandalone_rtio_core_sed_record15_payload_address2 = 2'd0;
reg [31:0] main_genericstandalone_rtio_core_sed_record15_payload_data2 = 32'd0;
reg main_genericstandalone_rtio_core_sed_replace_occured_r0 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r0 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory0_adr;
wire main_genericstandalone_rtio_core_sed_memory0_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r1 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r1 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory1_adr;
wire main_genericstandalone_rtio_core_sed_memory1_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r2 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r2 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory2_adr;
wire main_genericstandalone_rtio_core_sed_memory2_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r3 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r3 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory3_adr;
wire main_genericstandalone_rtio_core_sed_memory3_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r4 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r4 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory4_adr;
wire main_genericstandalone_rtio_core_sed_memory4_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r5 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r5 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory5_adr;
wire main_genericstandalone_rtio_core_sed_memory5_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r6 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r6 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory6_adr;
wire main_genericstandalone_rtio_core_sed_memory6_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r7 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r7 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory7_adr;
wire main_genericstandalone_rtio_core_sed_memory7_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r8 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r8 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory8_adr;
wire main_genericstandalone_rtio_core_sed_memory8_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r9 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r9 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory9_adr;
wire main_genericstandalone_rtio_core_sed_memory9_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r10 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r10 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory10_adr;
wire main_genericstandalone_rtio_core_sed_memory10_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r11 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r11 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory11_adr;
wire main_genericstandalone_rtio_core_sed_memory11_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r12 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r12 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory12_adr;
wire main_genericstandalone_rtio_core_sed_memory12_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r13 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r13 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory13_adr;
wire main_genericstandalone_rtio_core_sed_memory13_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r14 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r14 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory14_adr;
wire main_genericstandalone_rtio_core_sed_memory14_dat_r;
reg main_genericstandalone_rtio_core_sed_replace_occured_r15 = 1'd0;
reg main_genericstandalone_rtio_core_sed_nondata_replace_occured_r15 = 1'd0;
wire [5:0] main_genericstandalone_rtio_core_sed_memory15_adr;
wire main_genericstandalone_rtio_core_sed_memory15_dat_r;
wire main_genericstandalone_rtio_core_sed_selected0;
wire main_genericstandalone_rtio_core_sed_selected1;
wire main_genericstandalone_rtio_core_sed_selected2;
wire main_genericstandalone_rtio_core_sed_selected3;
wire main_genericstandalone_rtio_core_sed_selected4;
wire main_genericstandalone_rtio_core_sed_selected5;
wire main_genericstandalone_rtio_core_sed_selected6;
wire main_genericstandalone_rtio_core_sed_selected7;
wire main_genericstandalone_rtio_core_sed_selected8;
wire main_genericstandalone_rtio_core_sed_selected9;
wire main_genericstandalone_rtio_core_sed_selected10;
wire main_genericstandalone_rtio_core_sed_selected11;
wire main_genericstandalone_rtio_core_sed_selected12;
wire main_genericstandalone_rtio_core_sed_selected13;
wire main_genericstandalone_rtio_core_sed_selected14;
wire main_genericstandalone_rtio_core_sed_selected15;
wire main_genericstandalone_rtio_core_sed_selected16;
wire main_genericstandalone_rtio_core_sed_selected17;
wire main_genericstandalone_rtio_core_sed_selected18;
wire main_genericstandalone_rtio_core_sed_selected19;
wire main_genericstandalone_rtio_core_sed_selected20;
wire main_genericstandalone_rtio_core_sed_selected21;
wire main_genericstandalone_rtio_core_sed_selected22;
wire main_genericstandalone_rtio_core_sed_selected23;
wire main_genericstandalone_rtio_core_sed_selected24;
wire main_genericstandalone_rtio_core_sed_selected25;
wire main_genericstandalone_rtio_core_sed_selected26;
wire main_genericstandalone_rtio_core_sed_selected27;
wire main_genericstandalone_rtio_core_sed_selected28;
wire main_genericstandalone_rtio_core_sed_selected29;
wire main_genericstandalone_rtio_core_sed_selected30;
wire main_genericstandalone_rtio_core_sed_selected31;
wire main_genericstandalone_rtio_core_sed_selected32;
wire main_genericstandalone_rtio_core_sed_selected33;
wire main_genericstandalone_rtio_core_sed_selected34;
wire main_genericstandalone_rtio_core_sed_selected35;
wire main_genericstandalone_rtio_core_sed_selected36;
wire main_genericstandalone_rtio_core_sed_selected37;
wire main_genericstandalone_rtio_core_sed_selected38;
wire main_genericstandalone_rtio_core_sed_selected39;
wire main_genericstandalone_rtio_core_sed_selected40;
wire main_genericstandalone_rtio_core_sed_selected41;
wire main_genericstandalone_rtio_core_sed_selected42;
wire main_genericstandalone_rtio_core_sed_selected43;
wire main_genericstandalone_rtio_core_sed_selected44;
wire main_genericstandalone_rtio_core_sed_selected45;
wire main_genericstandalone_rtio_core_sed_selected46;
wire main_genericstandalone_rtio_core_sed_selected47;
wire main_genericstandalone_rtio_core_sed_selected48;
wire main_genericstandalone_rtio_core_sed_selected49;
wire main_genericstandalone_rtio_core_sed_selected50;
wire main_genericstandalone_rtio_core_sed_selected51;
wire main_genericstandalone_rtio_core_sed_selected52;
wire main_genericstandalone_rtio_core_sed_selected53;
wire main_genericstandalone_rtio_core_sed_selected54;
wire main_genericstandalone_rtio_core_sed_selected55;
wire main_genericstandalone_rtio_core_sed_selected56;
wire main_genericstandalone_rtio_core_sed_selected57;
wire main_genericstandalone_rtio_core_sed_selected58;
wire main_genericstandalone_rtio_core_sed_selected59;
wire main_genericstandalone_rtio_core_sed_selected60;
wire main_genericstandalone_rtio_core_sed_selected61;
wire main_genericstandalone_rtio_core_sed_selected62;
wire main_genericstandalone_rtio_core_sed_selected63;
wire main_genericstandalone_rtio_core_sed_selected64;
wire main_genericstandalone_rtio_core_sed_selected65;
wire main_genericstandalone_rtio_core_sed_selected66;
wire main_genericstandalone_rtio_core_sed_selected67;
wire main_genericstandalone_rtio_core_sed_selected68;
wire main_genericstandalone_rtio_core_sed_selected69;
wire main_genericstandalone_rtio_core_sed_selected70;
wire main_genericstandalone_rtio_core_sed_selected71;
wire main_genericstandalone_rtio_core_sed_selected72;
wire main_genericstandalone_rtio_core_sed_selected73;
wire main_genericstandalone_rtio_core_sed_selected74;
wire main_genericstandalone_rtio_core_sed_selected75;
wire main_genericstandalone_rtio_core_sed_selected76;
wire main_genericstandalone_rtio_core_sed_selected77;
wire main_genericstandalone_rtio_core_sed_selected78;
wire main_genericstandalone_rtio_core_sed_selected79;
wire main_genericstandalone_rtio_core_sed_selected80;
wire main_genericstandalone_rtio_core_sed_selected81;
wire main_genericstandalone_rtio_core_sed_selected82;
wire main_genericstandalone_rtio_core_sed_selected83;
wire main_genericstandalone_rtio_core_sed_selected84;
wire main_genericstandalone_rtio_core_sed_selected85;
wire main_genericstandalone_rtio_core_sed_selected86;
wire main_genericstandalone_rtio_core_sed_selected87;
wire main_genericstandalone_rtio_core_sed_selected88;
wire main_genericstandalone_rtio_core_sed_selected89;
wire main_genericstandalone_rtio_core_sed_selected90;
wire main_genericstandalone_rtio_core_sed_selected91;
wire main_genericstandalone_rtio_core_sed_selected92;
wire main_genericstandalone_rtio_core_sed_selected93;
wire main_genericstandalone_rtio_core_sed_selected94;
wire main_genericstandalone_rtio_core_sed_selected95;
wire main_genericstandalone_rtio_core_sed_selected96;
wire main_genericstandalone_rtio_core_sed_selected97;
wire main_genericstandalone_rtio_core_sed_selected98;
wire main_genericstandalone_rtio_core_sed_selected99;
wire main_genericstandalone_rtio_core_sed_selected100;
wire main_genericstandalone_rtio_core_sed_selected101;
wire main_genericstandalone_rtio_core_sed_selected102;
wire main_genericstandalone_rtio_core_sed_selected103;
wire main_genericstandalone_rtio_core_sed_selected104;
wire main_genericstandalone_rtio_core_sed_selected105;
wire main_genericstandalone_rtio_core_sed_selected106;
wire main_genericstandalone_rtio_core_sed_selected107;
wire main_genericstandalone_rtio_core_sed_selected108;
wire main_genericstandalone_rtio_core_sed_selected109;
wire main_genericstandalone_rtio_core_sed_selected110;
wire main_genericstandalone_rtio_core_sed_selected111;
wire main_genericstandalone_rtio_core_sed_selected112;
wire main_genericstandalone_rtio_core_sed_selected113;
wire main_genericstandalone_rtio_core_sed_selected114;
wire main_genericstandalone_rtio_core_sed_selected115;
wire main_genericstandalone_rtio_core_sed_selected116;
wire main_genericstandalone_rtio_core_sed_selected117;
wire main_genericstandalone_rtio_core_sed_selected118;
wire main_genericstandalone_rtio_core_sed_selected119;
wire main_genericstandalone_rtio_core_sed_selected120;
wire main_genericstandalone_rtio_core_sed_selected121;
wire main_genericstandalone_rtio_core_sed_selected122;
wire main_genericstandalone_rtio_core_sed_selected123;
wire main_genericstandalone_rtio_core_sed_selected124;
wire main_genericstandalone_rtio_core_sed_selected125;
wire main_genericstandalone_rtio_core_sed_selected126;
wire main_genericstandalone_rtio_core_sed_selected127;
wire main_genericstandalone_rtio_core_sed_selected128;
wire main_genericstandalone_rtio_core_sed_selected129;
wire main_genericstandalone_rtio_core_sed_selected130;
wire main_genericstandalone_rtio_core_sed_selected131;
wire main_genericstandalone_rtio_core_sed_selected132;
wire main_genericstandalone_rtio_core_sed_selected133;
wire main_genericstandalone_rtio_core_sed_selected134;
wire main_genericstandalone_rtio_core_sed_selected135;
wire main_genericstandalone_rtio_core_sed_selected136;
wire main_genericstandalone_rtio_core_sed_selected137;
wire main_genericstandalone_rtio_core_sed_selected138;
wire main_genericstandalone_rtio_core_sed_selected139;
wire main_genericstandalone_rtio_core_sed_selected140;
wire main_genericstandalone_rtio_core_sed_selected141;
wire main_genericstandalone_rtio_core_sed_selected142;
wire main_genericstandalone_rtio_core_sed_selected143;
wire main_genericstandalone_rtio_core_sed_selected144;
wire main_genericstandalone_rtio_core_sed_selected145;
wire main_genericstandalone_rtio_core_sed_selected146;
wire main_genericstandalone_rtio_core_sed_selected147;
wire main_genericstandalone_rtio_core_sed_selected148;
wire main_genericstandalone_rtio_core_sed_selected149;
wire main_genericstandalone_rtio_core_sed_selected150;
wire main_genericstandalone_rtio_core_sed_selected151;
wire main_genericstandalone_rtio_core_sed_selected152;
wire main_genericstandalone_rtio_core_sed_selected153;
wire main_genericstandalone_rtio_core_sed_selected154;
wire main_genericstandalone_rtio_core_sed_selected155;
wire main_genericstandalone_rtio_core_sed_selected156;
wire main_genericstandalone_rtio_core_sed_selected157;
wire main_genericstandalone_rtio_core_sed_selected158;
wire main_genericstandalone_rtio_core_sed_selected159;
wire main_genericstandalone_rtio_core_sed_selected160;
wire main_genericstandalone_rtio_core_sed_selected161;
wire main_genericstandalone_rtio_core_sed_selected162;
wire main_genericstandalone_rtio_core_sed_selected163;
wire main_genericstandalone_rtio_core_sed_selected164;
wire main_genericstandalone_rtio_core_sed_selected165;
wire main_genericstandalone_rtio_core_sed_selected166;
wire main_genericstandalone_rtio_core_sed_selected167;
wire main_genericstandalone_rtio_core_sed_selected168;
wire main_genericstandalone_rtio_core_sed_selected169;
wire main_genericstandalone_rtio_core_sed_selected170;
wire main_genericstandalone_rtio_core_sed_selected171;
wire main_genericstandalone_rtio_core_sed_selected172;
wire main_genericstandalone_rtio_core_sed_selected173;
wire main_genericstandalone_rtio_core_sed_selected174;
wire main_genericstandalone_rtio_core_sed_selected175;
wire main_genericstandalone_rtio_core_sed_selected176;
wire main_genericstandalone_rtio_core_sed_selected177;
wire main_genericstandalone_rtio_core_sed_selected178;
wire main_genericstandalone_rtio_core_sed_selected179;
wire main_genericstandalone_rtio_core_sed_selected180;
wire main_genericstandalone_rtio_core_sed_selected181;
wire main_genericstandalone_rtio_core_sed_selected182;
wire main_genericstandalone_rtio_core_sed_selected183;
wire main_genericstandalone_rtio_core_sed_selected184;
wire main_genericstandalone_rtio_core_sed_selected185;
wire main_genericstandalone_rtio_core_sed_selected186;
wire main_genericstandalone_rtio_core_sed_selected187;
wire main_genericstandalone_rtio_core_sed_selected188;
wire main_genericstandalone_rtio_core_sed_selected189;
wire main_genericstandalone_rtio_core_sed_selected190;
wire main_genericstandalone_rtio_core_sed_selected191;
wire main_genericstandalone_rtio_core_sed_selected192;
wire main_genericstandalone_rtio_core_sed_selected193;
wire main_genericstandalone_rtio_core_sed_selected194;
wire main_genericstandalone_rtio_core_sed_selected195;
wire main_genericstandalone_rtio_core_sed_selected196;
wire main_genericstandalone_rtio_core_sed_selected197;
wire main_genericstandalone_rtio_core_sed_selected198;
wire main_genericstandalone_rtio_core_sed_selected199;
wire main_genericstandalone_rtio_core_sed_selected200;
wire main_genericstandalone_rtio_core_sed_selected201;
wire main_genericstandalone_rtio_core_sed_selected202;
wire main_genericstandalone_rtio_core_sed_selected203;
wire main_genericstandalone_rtio_core_sed_selected204;
wire main_genericstandalone_rtio_core_sed_selected205;
wire main_genericstandalone_rtio_core_sed_selected206;
wire main_genericstandalone_rtio_core_sed_selected207;
wire main_genericstandalone_rtio_core_sed_selected208;
wire main_genericstandalone_rtio_core_sed_selected209;
wire main_genericstandalone_rtio_core_sed_selected210;
wire main_genericstandalone_rtio_core_sed_selected211;
wire main_genericstandalone_rtio_core_sed_selected212;
wire main_genericstandalone_rtio_core_sed_selected213;
wire main_genericstandalone_rtio_core_sed_selected214;
wire main_genericstandalone_rtio_core_sed_selected215;
wire main_genericstandalone_rtio_core_sed_selected216;
wire main_genericstandalone_rtio_core_sed_selected217;
wire main_genericstandalone_rtio_core_sed_selected218;
wire main_genericstandalone_rtio_core_sed_selected219;
wire main_genericstandalone_rtio_core_sed_selected220;
wire main_genericstandalone_rtio_core_sed_selected221;
wire main_genericstandalone_rtio_core_sed_selected222;
wire main_genericstandalone_rtio_core_sed_selected223;
wire main_genericstandalone_rtio_core_sed_selected224;
wire main_genericstandalone_rtio_core_sed_selected225;
wire main_genericstandalone_rtio_core_sed_selected226;
wire main_genericstandalone_rtio_core_sed_selected227;
wire main_genericstandalone_rtio_core_sed_selected228;
wire main_genericstandalone_rtio_core_sed_selected229;
wire main_genericstandalone_rtio_core_sed_selected230;
wire main_genericstandalone_rtio_core_sed_selected231;
wire main_genericstandalone_rtio_core_sed_selected232;
wire main_genericstandalone_rtio_core_sed_selected233;
wire main_genericstandalone_rtio_core_sed_selected234;
wire main_genericstandalone_rtio_core_sed_selected235;
wire main_genericstandalone_rtio_core_sed_selected236;
wire main_genericstandalone_rtio_core_sed_selected237;
wire main_genericstandalone_rtio_core_sed_selected238;
wire main_genericstandalone_rtio_core_sed_selected239;
wire main_genericstandalone_rtio_core_sed_selected240;
wire main_genericstandalone_rtio_core_sed_selected241;
wire main_genericstandalone_rtio_core_sed_selected242;
wire main_genericstandalone_rtio_core_sed_selected243;
wire main_genericstandalone_rtio_core_sed_selected244;
wire main_genericstandalone_rtio_core_sed_selected245;
wire main_genericstandalone_rtio_core_sed_selected246;
wire main_genericstandalone_rtio_core_sed_selected247;
wire main_genericstandalone_rtio_core_sed_selected248;
wire main_genericstandalone_rtio_core_sed_selected249;
wire main_genericstandalone_rtio_core_sed_selected250;
wire main_genericstandalone_rtio_core_sed_selected251;
wire main_genericstandalone_rtio_core_sed_selected252;
wire main_genericstandalone_rtio_core_sed_selected253;
wire main_genericstandalone_rtio_core_sed_selected254;
wire main_genericstandalone_rtio_core_sed_selected255;
wire main_genericstandalone_rtio_core_sed_selected256;
wire main_genericstandalone_rtio_core_sed_selected257;
wire main_genericstandalone_rtio_core_sed_selected258;
wire main_genericstandalone_rtio_core_sed_selected259;
wire main_genericstandalone_rtio_core_sed_selected260;
wire main_genericstandalone_rtio_core_sed_selected261;
wire main_genericstandalone_rtio_core_sed_selected262;
wire main_genericstandalone_rtio_core_sed_selected263;
wire main_genericstandalone_rtio_core_sed_selected264;
wire main_genericstandalone_rtio_core_sed_selected265;
wire main_genericstandalone_rtio_core_sed_selected266;
wire main_genericstandalone_rtio_core_sed_selected267;
wire main_genericstandalone_rtio_core_sed_selected268;
wire main_genericstandalone_rtio_core_sed_selected269;
wire main_genericstandalone_rtio_core_sed_selected270;
wire main_genericstandalone_rtio_core_sed_selected271;
wire main_genericstandalone_rtio_core_sed_selected272;
wire main_genericstandalone_rtio_core_sed_selected273;
wire main_genericstandalone_rtio_core_sed_selected274;
wire main_genericstandalone_rtio_core_sed_selected275;
wire main_genericstandalone_rtio_core_sed_selected276;
wire main_genericstandalone_rtio_core_sed_selected277;
wire main_genericstandalone_rtio_core_sed_selected278;
wire main_genericstandalone_rtio_core_sed_selected279;
wire main_genericstandalone_rtio_core_sed_selected280;
wire main_genericstandalone_rtio_core_sed_selected281;
wire main_genericstandalone_rtio_core_sed_selected282;
wire main_genericstandalone_rtio_core_sed_selected283;
wire main_genericstandalone_rtio_core_sed_selected284;
wire main_genericstandalone_rtio_core_sed_selected285;
wire main_genericstandalone_rtio_core_sed_selected286;
wire main_genericstandalone_rtio_core_sed_selected287;
wire main_genericstandalone_rtio_core_sed_selected288;
wire main_genericstandalone_rtio_core_sed_selected289;
wire main_genericstandalone_rtio_core_sed_selected290;
wire main_genericstandalone_rtio_core_sed_selected291;
wire main_genericstandalone_rtio_core_sed_selected292;
wire main_genericstandalone_rtio_core_sed_selected293;
wire main_genericstandalone_rtio_core_sed_selected294;
wire main_genericstandalone_rtio_core_sed_selected295;
wire main_genericstandalone_rtio_core_sed_selected296;
wire main_genericstandalone_rtio_core_sed_selected297;
wire main_genericstandalone_rtio_core_sed_selected298;
wire main_genericstandalone_rtio_core_sed_selected299;
wire main_genericstandalone_rtio_core_sed_selected300;
wire main_genericstandalone_rtio_core_sed_selected301;
wire main_genericstandalone_rtio_core_sed_selected302;
wire main_genericstandalone_rtio_core_sed_selected303;
wire main_genericstandalone_rtio_core_sed_selected304;
wire main_genericstandalone_rtio_core_sed_selected305;
wire main_genericstandalone_rtio_core_sed_selected306;
wire main_genericstandalone_rtio_core_sed_selected307;
wire main_genericstandalone_rtio_core_sed_selected308;
wire main_genericstandalone_rtio_core_sed_selected309;
wire main_genericstandalone_rtio_core_sed_selected310;
wire main_genericstandalone_rtio_core_sed_selected311;
wire main_genericstandalone_rtio_core_sed_selected312;
wire main_genericstandalone_rtio_core_sed_selected313;
wire main_genericstandalone_rtio_core_sed_selected314;
wire main_genericstandalone_rtio_core_sed_selected315;
wire main_genericstandalone_rtio_core_sed_selected316;
wire main_genericstandalone_rtio_core_sed_selected317;
wire main_genericstandalone_rtio_core_sed_selected318;
wire main_genericstandalone_rtio_core_sed_selected319;
wire main_genericstandalone_rtio_core_sed_selected320;
wire main_genericstandalone_rtio_core_sed_selected321;
wire main_genericstandalone_rtio_core_sed_selected322;
wire main_genericstandalone_rtio_core_sed_selected323;
wire main_genericstandalone_rtio_core_sed_selected324;
wire main_genericstandalone_rtio_core_sed_selected325;
wire main_genericstandalone_rtio_core_sed_selected326;
wire main_genericstandalone_rtio_core_sed_selected327;
wire main_genericstandalone_rtio_core_sed_selected328;
wire main_genericstandalone_rtio_core_sed_selected329;
wire main_genericstandalone_rtio_core_sed_selected330;
wire main_genericstandalone_rtio_core_sed_selected331;
wire main_genericstandalone_rtio_core_sed_selected332;
wire main_genericstandalone_rtio_core_sed_selected333;
wire main_genericstandalone_rtio_core_sed_selected334;
wire main_genericstandalone_rtio_core_sed_selected335;
wire main_genericstandalone_rtio_core_sed_selected336;
wire main_genericstandalone_rtio_core_sed_selected337;
wire main_genericstandalone_rtio_core_sed_selected338;
wire main_genericstandalone_rtio_core_sed_selected339;
wire main_genericstandalone_rtio_core_sed_selected340;
wire main_genericstandalone_rtio_core_sed_selected341;
wire main_genericstandalone_rtio_core_sed_selected342;
wire main_genericstandalone_rtio_core_sed_selected343;
wire main_genericstandalone_rtio_core_sed_selected344;
wire main_genericstandalone_rtio_core_sed_selected345;
wire main_genericstandalone_rtio_core_sed_selected346;
wire main_genericstandalone_rtio_core_sed_selected347;
wire main_genericstandalone_rtio_core_sed_selected348;
wire main_genericstandalone_rtio_core_sed_selected349;
wire main_genericstandalone_rtio_core_sed_selected350;
wire main_genericstandalone_rtio_core_sed_selected351;
wire main_genericstandalone_rtio_core_sed_selected352;
wire main_genericstandalone_rtio_core_sed_selected353;
wire main_genericstandalone_rtio_core_sed_selected354;
wire main_genericstandalone_rtio_core_sed_selected355;
wire main_genericstandalone_rtio_core_sed_selected356;
wire main_genericstandalone_rtio_core_sed_selected357;
wire main_genericstandalone_rtio_core_sed_selected358;
wire main_genericstandalone_rtio_core_sed_selected359;
wire main_genericstandalone_rtio_core_sed_selected360;
wire main_genericstandalone_rtio_core_sed_selected361;
wire main_genericstandalone_rtio_core_sed_selected362;
wire main_genericstandalone_rtio_core_sed_selected363;
wire main_genericstandalone_rtio_core_sed_selected364;
wire main_genericstandalone_rtio_core_sed_selected365;
wire main_genericstandalone_rtio_core_sed_selected366;
wire main_genericstandalone_rtio_core_sed_selected367;
wire main_genericstandalone_rtio_core_sed_selected368;
wire main_genericstandalone_rtio_core_sed_selected369;
wire main_genericstandalone_rtio_core_sed_selected370;
wire main_genericstandalone_rtio_core_sed_selected371;
wire main_genericstandalone_rtio_core_sed_selected372;
wire main_genericstandalone_rtio_core_sed_selected373;
wire main_genericstandalone_rtio_core_sed_selected374;
wire main_genericstandalone_rtio_core_sed_selected375;
wire main_genericstandalone_rtio_core_sed_selected376;
wire main_genericstandalone_rtio_core_sed_selected377;
wire main_genericstandalone_rtio_core_sed_selected378;
wire main_genericstandalone_rtio_core_sed_selected379;
wire main_genericstandalone_rtio_core_sed_selected380;
wire main_genericstandalone_rtio_core_sed_selected381;
wire main_genericstandalone_rtio_core_sed_selected382;
wire main_genericstandalone_rtio_core_sed_selected383;
wire main_genericstandalone_rtio_core_sed_selected384;
wire main_genericstandalone_rtio_core_sed_selected385;
wire main_genericstandalone_rtio_core_sed_selected386;
wire main_genericstandalone_rtio_core_sed_selected387;
wire main_genericstandalone_rtio_core_sed_selected388;
wire main_genericstandalone_rtio_core_sed_selected389;
wire main_genericstandalone_rtio_core_sed_selected390;
wire main_genericstandalone_rtio_core_sed_selected391;
wire main_genericstandalone_rtio_core_sed_selected392;
wire main_genericstandalone_rtio_core_sed_selected393;
wire main_genericstandalone_rtio_core_sed_selected394;
wire main_genericstandalone_rtio_core_sed_selected395;
wire main_genericstandalone_rtio_core_sed_selected396;
wire main_genericstandalone_rtio_core_sed_selected397;
wire main_genericstandalone_rtio_core_sed_selected398;
wire main_genericstandalone_rtio_core_sed_selected399;
wire main_genericstandalone_rtio_core_sed_selected400;
wire main_genericstandalone_rtio_core_sed_selected401;
wire main_genericstandalone_rtio_core_sed_selected402;
wire main_genericstandalone_rtio_core_sed_selected403;
wire main_genericstandalone_rtio_core_sed_selected404;
wire main_genericstandalone_rtio_core_sed_selected405;
wire main_genericstandalone_rtio_core_sed_selected406;
wire main_genericstandalone_rtio_core_sed_selected407;
wire main_genericstandalone_rtio_core_sed_selected408;
wire main_genericstandalone_rtio_core_sed_selected409;
wire main_genericstandalone_rtio_core_sed_selected410;
wire main_genericstandalone_rtio_core_sed_selected411;
wire main_genericstandalone_rtio_core_sed_selected412;
wire main_genericstandalone_rtio_core_sed_selected413;
wire main_genericstandalone_rtio_core_sed_selected414;
wire main_genericstandalone_rtio_core_sed_selected415;
wire main_genericstandalone_rtio_core_sed_selected416;
wire main_genericstandalone_rtio_core_sed_selected417;
wire main_genericstandalone_rtio_core_sed_selected418;
wire main_genericstandalone_rtio_core_sed_selected419;
wire main_genericstandalone_rtio_core_sed_selected420;
wire main_genericstandalone_rtio_core_sed_selected421;
wire main_genericstandalone_rtio_core_sed_selected422;
wire main_genericstandalone_rtio_core_sed_selected423;
wire main_genericstandalone_rtio_core_sed_selected424;
wire main_genericstandalone_rtio_core_sed_selected425;
wire main_genericstandalone_rtio_core_sed_selected426;
wire main_genericstandalone_rtio_core_sed_selected427;
wire main_genericstandalone_rtio_core_sed_selected428;
wire main_genericstandalone_rtio_core_sed_selected429;
wire main_genericstandalone_rtio_core_sed_selected430;
wire main_genericstandalone_rtio_core_sed_selected431;
wire main_genericstandalone_rtio_core_sed_selected432;
wire main_genericstandalone_rtio_core_sed_selected433;
wire main_genericstandalone_rtio_core_sed_selected434;
wire main_genericstandalone_rtio_core_sed_selected435;
wire main_genericstandalone_rtio_core_sed_selected436;
wire main_genericstandalone_rtio_core_sed_selected437;
wire main_genericstandalone_rtio_core_sed_selected438;
wire main_genericstandalone_rtio_core_sed_selected439;
wire main_genericstandalone_rtio_core_sed_selected440;
wire main_genericstandalone_rtio_core_sed_selected441;
wire main_genericstandalone_rtio_core_sed_selected442;
wire main_genericstandalone_rtio_core_sed_selected443;
wire main_genericstandalone_rtio_core_sed_selected444;
wire main_genericstandalone_rtio_core_sed_selected445;
wire main_genericstandalone_rtio_core_sed_selected446;
wire main_genericstandalone_rtio_core_sed_selected447;
wire main_genericstandalone_rtio_core_sed_selected448;
wire main_genericstandalone_rtio_core_sed_selected449;
wire main_genericstandalone_rtio_core_sed_selected450;
wire main_genericstandalone_rtio_core_sed_selected451;
wire main_genericstandalone_rtio_core_sed_selected452;
wire main_genericstandalone_rtio_core_sed_selected453;
wire main_genericstandalone_rtio_core_sed_selected454;
wire main_genericstandalone_rtio_core_sed_selected455;
wire main_genericstandalone_rtio_core_sed_selected456;
wire main_genericstandalone_rtio_core_sed_selected457;
wire main_genericstandalone_rtio_core_sed_selected458;
wire main_genericstandalone_rtio_core_sed_selected459;
wire main_genericstandalone_rtio_core_sed_selected460;
wire main_genericstandalone_rtio_core_sed_selected461;
wire main_genericstandalone_rtio_core_sed_selected462;
wire main_genericstandalone_rtio_core_sed_selected463;
wire main_genericstandalone_rtio_core_sed_selected464;
wire main_genericstandalone_rtio_core_sed_selected465;
wire main_genericstandalone_rtio_core_sed_selected466;
wire main_genericstandalone_rtio_core_sed_selected467;
wire main_genericstandalone_rtio_core_sed_selected468;
wire main_genericstandalone_rtio_core_sed_selected469;
wire main_genericstandalone_rtio_core_sed_selected470;
wire main_genericstandalone_rtio_core_sed_selected471;
wire main_genericstandalone_rtio_core_sed_selected472;
wire main_genericstandalone_rtio_core_sed_selected473;
wire main_genericstandalone_rtio_core_sed_selected474;
wire main_genericstandalone_rtio_core_sed_selected475;
wire main_genericstandalone_rtio_core_sed_selected476;
wire main_genericstandalone_rtio_core_sed_selected477;
wire main_genericstandalone_rtio_core_sed_selected478;
wire main_genericstandalone_rtio_core_sed_selected479;
wire main_genericstandalone_rtio_core_sed_selected480;
wire main_genericstandalone_rtio_core_sed_selected481;
wire main_genericstandalone_rtio_core_sed_selected482;
wire main_genericstandalone_rtio_core_sed_selected483;
wire main_genericstandalone_rtio_core_sed_selected484;
wire main_genericstandalone_rtio_core_sed_selected485;
wire main_genericstandalone_rtio_core_sed_selected486;
wire main_genericstandalone_rtio_core_sed_selected487;
wire main_genericstandalone_rtio_core_sed_selected488;
wire main_genericstandalone_rtio_core_sed_selected489;
wire main_genericstandalone_rtio_core_sed_selected490;
wire main_genericstandalone_rtio_core_sed_selected491;
wire main_genericstandalone_rtio_core_sed_selected492;
wire main_genericstandalone_rtio_core_sed_selected493;
wire main_genericstandalone_rtio_core_sed_selected494;
wire main_genericstandalone_rtio_core_sed_selected495;
wire main_genericstandalone_rtio_core_sed_selected496;
wire main_genericstandalone_rtio_core_sed_selected497;
wire main_genericstandalone_rtio_core_sed_selected498;
wire main_genericstandalone_rtio_core_sed_selected499;
wire main_genericstandalone_rtio_core_sed_selected500;
wire main_genericstandalone_rtio_core_sed_selected501;
wire main_genericstandalone_rtio_core_sed_selected502;
wire main_genericstandalone_rtio_core_sed_selected503;
wire main_genericstandalone_rtio_core_sed_selected504;
wire main_genericstandalone_rtio_core_sed_selected505;
wire main_genericstandalone_rtio_core_sed_selected506;
wire main_genericstandalone_rtio_core_sed_selected507;
wire main_genericstandalone_rtio_core_sed_selected508;
wire main_genericstandalone_rtio_core_sed_selected509;
wire main_genericstandalone_rtio_core_sed_selected510;
wire main_genericstandalone_rtio_core_sed_selected511;
wire main_genericstandalone_rtio_core_sed_selected512;
wire main_genericstandalone_rtio_core_sed_selected513;
wire main_genericstandalone_rtio_core_sed_selected514;
wire main_genericstandalone_rtio_core_sed_selected515;
wire main_genericstandalone_rtio_core_sed_selected516;
wire main_genericstandalone_rtio_core_sed_selected517;
wire main_genericstandalone_rtio_core_sed_selected518;
wire main_genericstandalone_rtio_core_sed_selected519;
wire main_genericstandalone_rtio_core_sed_selected520;
wire main_genericstandalone_rtio_core_sed_selected521;
wire main_genericstandalone_rtio_core_sed_selected522;
wire main_genericstandalone_rtio_core_sed_selected523;
wire main_genericstandalone_rtio_core_sed_selected524;
wire main_genericstandalone_rtio_core_sed_selected525;
wire main_genericstandalone_rtio_core_sed_selected526;
wire main_genericstandalone_rtio_core_sed_selected527;
wire main_genericstandalone_rtio_core_sed_selected528;
wire main_genericstandalone_rtio_core_sed_selected529;
wire main_genericstandalone_rtio_core_sed_selected530;
wire main_genericstandalone_rtio_core_sed_selected531;
wire main_genericstandalone_rtio_core_sed_selected532;
wire main_genericstandalone_rtio_core_sed_selected533;
wire main_genericstandalone_rtio_core_sed_selected534;
wire main_genericstandalone_rtio_core_sed_selected535;
wire main_genericstandalone_rtio_core_sed_selected536;
wire main_genericstandalone_rtio_core_sed_selected537;
wire main_genericstandalone_rtio_core_sed_selected538;
wire main_genericstandalone_rtio_core_sed_selected539;
wire main_genericstandalone_rtio_core_sed_selected540;
wire main_genericstandalone_rtio_core_sed_selected541;
wire main_genericstandalone_rtio_core_sed_selected542;
wire main_genericstandalone_rtio_core_sed_selected543;
wire main_genericstandalone_rtio_core_sed_selected544;
wire main_genericstandalone_rtio_core_sed_selected545;
wire main_genericstandalone_rtio_core_sed_selected546;
wire main_genericstandalone_rtio_core_sed_selected547;
wire main_genericstandalone_rtio_core_sed_selected548;
wire main_genericstandalone_rtio_core_sed_selected549;
wire main_genericstandalone_rtio_core_sed_selected550;
wire main_genericstandalone_rtio_core_sed_selected551;
wire main_genericstandalone_rtio_core_sed_selected552;
wire main_genericstandalone_rtio_core_sed_selected553;
wire main_genericstandalone_rtio_core_sed_selected554;
wire main_genericstandalone_rtio_core_sed_selected555;
wire main_genericstandalone_rtio_core_sed_selected556;
wire main_genericstandalone_rtio_core_sed_selected557;
wire main_genericstandalone_rtio_core_sed_selected558;
wire main_genericstandalone_rtio_core_sed_selected559;
wire main_genericstandalone_rtio_core_sed_selected560;
wire main_genericstandalone_rtio_core_sed_selected561;
wire main_genericstandalone_rtio_core_sed_selected562;
wire main_genericstandalone_rtio_core_sed_selected563;
wire main_genericstandalone_rtio_core_sed_selected564;
wire main_genericstandalone_rtio_core_sed_selected565;
wire main_genericstandalone_rtio_core_sed_selected566;
wire main_genericstandalone_rtio_core_sed_selected567;
wire main_genericstandalone_rtio_core_sed_selected568;
wire main_genericstandalone_rtio_core_sed_selected569;
wire main_genericstandalone_rtio_core_sed_selected570;
wire main_genericstandalone_rtio_core_sed_selected571;
wire main_genericstandalone_rtio_core_sed_selected572;
wire main_genericstandalone_rtio_core_sed_selected573;
wire main_genericstandalone_rtio_core_sed_selected574;
wire main_genericstandalone_rtio_core_sed_selected575;
wire main_genericstandalone_rtio_core_sed_selected576;
wire main_genericstandalone_rtio_core_sed_selected577;
wire main_genericstandalone_rtio_core_sed_selected578;
wire main_genericstandalone_rtio_core_sed_selected579;
wire main_genericstandalone_rtio_core_sed_selected580;
wire main_genericstandalone_rtio_core_sed_selected581;
wire main_genericstandalone_rtio_core_sed_selected582;
wire main_genericstandalone_rtio_core_sed_selected583;
wire main_genericstandalone_rtio_core_sed_selected584;
wire main_genericstandalone_rtio_core_sed_selected585;
wire main_genericstandalone_rtio_core_sed_selected586;
wire main_genericstandalone_rtio_core_sed_selected587;
wire main_genericstandalone_rtio_core_sed_selected588;
wire main_genericstandalone_rtio_core_sed_selected589;
wire main_genericstandalone_rtio_core_sed_selected590;
wire main_genericstandalone_rtio_core_sed_selected591;
wire main_genericstandalone_rtio_core_sed_selected592;
wire main_genericstandalone_rtio_core_sed_selected593;
wire main_genericstandalone_rtio_core_sed_selected594;
wire main_genericstandalone_rtio_core_sed_selected595;
wire main_genericstandalone_rtio_core_sed_selected596;
wire main_genericstandalone_rtio_core_sed_selected597;
wire main_genericstandalone_rtio_core_sed_selected598;
wire main_genericstandalone_rtio_core_sed_selected599;
wire main_genericstandalone_rtio_core_sed_selected600;
wire main_genericstandalone_rtio_core_sed_selected601;
wire main_genericstandalone_rtio_core_sed_selected602;
wire main_genericstandalone_rtio_core_sed_selected603;
wire main_genericstandalone_rtio_core_sed_selected604;
wire main_genericstandalone_rtio_core_sed_selected605;
wire main_genericstandalone_rtio_core_sed_selected606;
wire main_genericstandalone_rtio_core_sed_selected607;
reg main_genericstandalone_rtio_core_sed_stb_r0 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r0 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r1 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r1 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r2 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r2 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r3 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r3 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r4 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r4 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r5 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r5 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r6 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r6 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r7 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r7 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r8 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r8 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r9 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r9 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r10 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r10 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r11 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r11 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r12 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r12 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r13 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r13 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r14 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r14 = 6'd0;
reg main_genericstandalone_rtio_core_sed_stb_r15 = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_sed_channel_r15 = 6'd0;
reg main_genericstandalone_rtio_core_inputcollector_i_ack = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_readable;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_din;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_dout;
reg [6:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 = 7'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_replace = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_produce = 6'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_consume = 6'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_adr;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_we;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_do_read;
wire [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_adr;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_re;
wire [6:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level1;
wire main_genericstandalone_rtio_core_inputcollector_record0_fifo_in_data;
wire [63:0] main_genericstandalone_rtio_core_inputcollector_record0_fifo_in_timestamp;
wire main_genericstandalone_rtio_core_inputcollector_record0_fifo_out_data;
wire [63:0] main_genericstandalone_rtio_core_inputcollector_record0_fifo_out_timestamp;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger0;
wire main_genericstandalone_rtio_core_inputcollector_selected0;
reg main_genericstandalone_rtio_core_inputcollector_overflow0 = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_readable;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_din;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_dout;
reg [6:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 = 7'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_replace = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_produce = 6'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_consume = 6'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_adr;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_we;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_do_read;
wire [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_adr;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_re;
wire [6:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level1;
wire main_genericstandalone_rtio_core_inputcollector_record1_fifo_in_data;
wire [63:0] main_genericstandalone_rtio_core_inputcollector_record1_fifo_in_timestamp;
wire main_genericstandalone_rtio_core_inputcollector_record1_fifo_out_data;
wire [63:0] main_genericstandalone_rtio_core_inputcollector_record1_fifo_out_timestamp;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger1;
wire main_genericstandalone_rtio_core_inputcollector_selected1;
reg main_genericstandalone_rtio_core_inputcollector_overflow1 = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_readable;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_din;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_dout;
reg [6:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 = 7'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_replace = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_produce = 6'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_consume = 6'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_adr;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_we;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_do_read;
wire [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_adr;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_re;
wire [6:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level1;
wire main_genericstandalone_rtio_core_inputcollector_record2_fifo_in_data;
wire [63:0] main_genericstandalone_rtio_core_inputcollector_record2_fifo_in_timestamp;
wire main_genericstandalone_rtio_core_inputcollector_record2_fifo_out_data;
wire [63:0] main_genericstandalone_rtio_core_inputcollector_record2_fifo_out_timestamp;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger2;
wire main_genericstandalone_rtio_core_inputcollector_selected2;
reg main_genericstandalone_rtio_core_inputcollector_overflow2 = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_readable;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_din;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_dout;
reg [6:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 = 7'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_replace = 1'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_produce = 6'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_consume = 6'd0;
reg [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_adr;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_we;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_do_read;
wire [5:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_adr;
wire [64:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_re;
wire [6:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level1;
wire main_genericstandalone_rtio_core_inputcollector_record3_fifo_in_data;
wire [63:0] main_genericstandalone_rtio_core_inputcollector_record3_fifo_in_timestamp;
wire main_genericstandalone_rtio_core_inputcollector_record3_fifo_out_data;
wire [63:0] main_genericstandalone_rtio_core_inputcollector_record3_fifo_out_timestamp;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger3;
wire main_genericstandalone_rtio_core_inputcollector_selected3;
reg main_genericstandalone_rtio_core_inputcollector_overflow3 = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_readable;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_din;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_dout;
reg [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 = 3'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_replace = 1'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_produce = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_consume = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_we;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_do_read;
wire [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_re;
wire [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level1;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record4_fifo_in_data;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record4_fifo_out_data;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger4;
wire main_genericstandalone_rtio_core_inputcollector_selected4;
reg main_genericstandalone_rtio_core_inputcollector_overflow4 = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_readable;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_din;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_dout;
reg [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 = 3'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_replace = 1'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_produce = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_consume = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_we;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_do_read;
wire [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_re;
wire [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level1;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record5_fifo_in_data;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record5_fifo_out_data;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger5;
wire main_genericstandalone_rtio_core_inputcollector_selected5;
reg main_genericstandalone_rtio_core_inputcollector_overflow5 = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_readable;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_din;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_dout;
reg [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 = 3'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_replace = 1'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_produce = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_consume = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_we;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_do_read;
wire [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_re;
wire [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level1;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record6_fifo_in_data;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record6_fifo_out_data;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger6;
wire main_genericstandalone_rtio_core_inputcollector_selected6;
reg main_genericstandalone_rtio_core_inputcollector_overflow6 = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_readable;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_din;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_dout;
reg [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 = 3'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_replace = 1'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_produce = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_consume = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_we;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_do_read;
wire [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_re;
wire [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level1;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record7_fifo_in_data;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record7_fifo_out_data;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger7;
wire main_genericstandalone_rtio_core_inputcollector_selected7;
reg main_genericstandalone_rtio_core_inputcollector_overflow7 = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_re;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_readable = 1'd0;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_we;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_writable;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_re;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_readable;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_din;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_dout;
reg [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 = 3'd0;
reg main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_replace = 1'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_produce = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_consume = 2'd0;
reg [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_we;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_dat_w;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_do_read;
wire [1:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_adr;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_dat_r;
wire main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_re;
wire [2:0] main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level1;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record8_fifo_in_data;
wire [31:0] main_genericstandalone_rtio_core_inputcollector_record8_fifo_out_data;
wire main_genericstandalone_rtio_core_inputcollector_overflow_trigger8;
wire main_genericstandalone_rtio_core_inputcollector_selected8;
reg main_genericstandalone_rtio_core_inputcollector_overflow8 = 1'd0;
wire [1:0] main_genericstandalone_rtio_core_inputcollector_i_status_raw;
reg [63:0] main_genericstandalone_rtio_core_inputcollector_input_timeout = 64'd0;
reg main_genericstandalone_rtio_core_inputcollector_input_pending = 1'd0;
wire main_genericstandalone_rtio_core_o_collision_sync_i;
wire main_genericstandalone_rtio_core_o_collision_sync_o;
wire [15:0] main_genericstandalone_rtio_core_o_collision_sync_data_i;
wire [15:0] main_genericstandalone_rtio_core_o_collision_sync_data_o;
wire main_genericstandalone_rtio_core_o_collision_sync_ps_i;
wire main_genericstandalone_rtio_core_o_collision_sync_ps_o;
reg main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_i = 1'd0;
wire main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_o;
reg main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_o_r = 1'd0;
wire main_genericstandalone_rtio_core_o_collision_sync_ps_ack_i;
wire main_genericstandalone_rtio_core_o_collision_sync_ps_ack_o;
reg main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_i = 1'd0;
wire main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_o;
reg main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_o_r = 1'd0;
reg main_genericstandalone_rtio_core_o_collision_sync_blind = 1'd0;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_rtio_core_o_collision_sync_bxfer_data = 16'd0;
wire main_genericstandalone_rtio_core_o_busy_sync_i;
wire main_genericstandalone_rtio_core_o_busy_sync_o;
wire [15:0] main_genericstandalone_rtio_core_o_busy_sync_data_i;
wire [15:0] main_genericstandalone_rtio_core_o_busy_sync_data_o;
wire main_genericstandalone_rtio_core_o_busy_sync_ps_i;
wire main_genericstandalone_rtio_core_o_busy_sync_ps_o;
reg main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_i = 1'd0;
wire main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_o;
reg main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_o_r = 1'd0;
wire main_genericstandalone_rtio_core_o_busy_sync_ps_ack_i;
wire main_genericstandalone_rtio_core_o_busy_sync_ps_ack_o;
reg main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_i = 1'd0;
wire main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_o;
reg main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_o_r = 1'd0;
reg main_genericstandalone_rtio_core_o_busy_sync_blind = 1'd0;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_rtio_core_o_busy_sync_bxfer_data = 16'd0;
reg main_genericstandalone_rtio_core_o_collision = 1'd0;
reg main_genericstandalone_rtio_core_o_busy = 1'd0;
reg main_genericstandalone_rtio_core_o_sequence_error = 1'd0;
reg [31:0] main_genericstandalone_rtio_target_storage_full = 32'd0;
wire [31:0] main_genericstandalone_rtio_target_storage;
reg main_genericstandalone_rtio_target_re = 1'd0;
wire main_genericstandalone_rtio_now_hi_re;
wire [31:0] main_genericstandalone_rtio_now_hi_r;
wire [31:0] main_genericstandalone_rtio_now_hi_w;
wire main_genericstandalone_rtio_now_lo_re;
wire [31:0] main_genericstandalone_rtio_now_lo_r;
wire [31:0] main_genericstandalone_rtio_now_lo_w;
reg [511:0] main_genericstandalone_rtio_o_data_storage_full = 512'd0;
wire [511:0] main_genericstandalone_rtio_o_data_storage;
reg main_genericstandalone_rtio_o_data_re = 1'd0;
wire main_genericstandalone_rtio_o_data_we;
wire [511:0] main_genericstandalone_rtio_o_data_dat_w;
wire [2:0] main_genericstandalone_rtio_o_status_status;
reg [63:0] main_genericstandalone_rtio_i_timeout_storage_full = 64'd0;
wire [63:0] main_genericstandalone_rtio_i_timeout_storage;
reg main_genericstandalone_rtio_i_timeout_re = 1'd0;
wire [31:0] main_genericstandalone_rtio_i_data_status;
wire [63:0] main_genericstandalone_rtio_i_timestamp_status;
wire [3:0] main_genericstandalone_rtio_i_status_status;
reg [63:0] main_genericstandalone_rtio_counter_status = 64'd0;
wire main_genericstandalone_rtio_counter_update_re;
wire main_genericstandalone_rtio_counter_update_r;
reg main_genericstandalone_rtio_counter_update_w = 1'd0;
reg [1:0] main_genericstandalone_rtio_cri_cmd;
wire [23:0] main_genericstandalone_rtio_cri_chan_sel;
wire [63:0] main_genericstandalone_rtio_cri_o_timestamp;
wire [511:0] main_genericstandalone_rtio_cri_o_data;
wire [7:0] main_genericstandalone_rtio_cri_o_address;
wire [2:0] main_genericstandalone_rtio_cri_o_status;
wire main_genericstandalone_rtio_cri_o_buffer_space_valid;
wire [15:0] main_genericstandalone_rtio_cri_o_buffer_space;
wire [63:0] main_genericstandalone_rtio_cri_i_timeout;
wire [31:0] main_genericstandalone_rtio_cri_i_data;
wire [63:0] main_genericstandalone_rtio_cri_i_timestamp;
wire [3:0] main_genericstandalone_rtio_cri_i_status;
reg [63:0] main_genericstandalone_rtio_now = 64'd0;
reg [31:0] main_genericstandalone_rtio_now_hi_backing = 32'd0;
wire [28:0] main_genericstandalone_interface0_bus_adr;
reg [127:0] main_genericstandalone_interface0_bus_dat_w = 128'd0;
wire [127:0] main_genericstandalone_interface0_bus_dat_r;
reg [15:0] main_genericstandalone_interface0_bus_sel = 16'd0;
wire main_genericstandalone_interface0_bus_cyc;
wire main_genericstandalone_interface0_bus_stb;
wire main_genericstandalone_interface0_bus_ack;
reg main_genericstandalone_interface0_bus_we = 1'd0;
wire [2:0] main_genericstandalone_interface0_bus_cti;
reg [1:0] main_genericstandalone_interface0_bus_bte = 2'd0;
wire main_genericstandalone_interface0_bus_err;
wire main_genericstandalone_dma_enable_enable_re;
wire main_genericstandalone_dma_enable_enable_r;
reg main_genericstandalone_dma_enable_enable_w;
reg main_genericstandalone_dma_flow_enable;
reg main_genericstandalone_dma_dma_sink_stb = 1'd0;
wire main_genericstandalone_dma_dma_sink_ack;
reg main_genericstandalone_dma_dma_sink_eop = 1'd0;
reg [28:0] main_genericstandalone_dma_dma_sink_payload_address = 29'd0;
wire main_genericstandalone_dma_dma_source_stb;
wire main_genericstandalone_dma_dma_source_ack;
wire main_genericstandalone_dma_dma_source_last;
wire main_genericstandalone_dma_dma_source_eop;
wire [127:0] main_genericstandalone_dma_dma_source_payload_data;
wire main_genericstandalone_dma_dma_bus_stb;
reg [5:0] main_genericstandalone_dma_dma_transfer_cyc = 6'd63;
wire main_genericstandalone_dma_dma_transfer_cyc_ce;
wire main_genericstandalone_dma_dma_transfer_cyc_rst;
wire main_genericstandalone_dma_dma_last;
reg [32:0] main_genericstandalone_dma_dma_storage_full = 33'd0;
wire [28:0] main_genericstandalone_dma_dma_storage;
reg main_genericstandalone_dma_dma_re = 1'd0;
reg main_genericstandalone_dma_dma_enable_r = 1'd0;
wire main_genericstandalone_dma_fifo_sink_stb;
reg main_genericstandalone_dma_fifo_sink_ack;
wire main_genericstandalone_dma_fifo_sink_last;
wire main_genericstandalone_dma_fifo_sink_eop;
wire [127:0] main_genericstandalone_dma_fifo_sink_payload_data;
wire main_genericstandalone_dma_fifo_source_stb;
wire main_genericstandalone_dma_fifo_source_ack;
reg main_genericstandalone_dma_fifo_source_last = 1'd0;
wire main_genericstandalone_dma_fifo_source_eop;
wire [127:0] main_genericstandalone_dma_fifo_source_payload_data;
wire main_genericstandalone_dma_fifo_re;
reg main_genericstandalone_dma_fifo_readable = 1'd0;
reg main_genericstandalone_dma_fifo_syncfifo_we;
wire main_genericstandalone_dma_fifo_syncfifo_writable;
wire main_genericstandalone_dma_fifo_syncfifo_re;
wire main_genericstandalone_dma_fifo_syncfifo_readable;
wire [128:0] main_genericstandalone_dma_fifo_syncfifo_din;
wire [128:0] main_genericstandalone_dma_fifo_syncfifo_dout;
reg [7:0] main_genericstandalone_dma_fifo_level0 = 8'd0;
reg main_genericstandalone_dma_fifo_replace = 1'd0;
reg [6:0] main_genericstandalone_dma_fifo_produce = 7'd0;
reg [6:0] main_genericstandalone_dma_fifo_consume = 7'd0;
reg [6:0] main_genericstandalone_dma_fifo_wrport_adr;
wire [128:0] main_genericstandalone_dma_fifo_wrport_dat_r;
wire main_genericstandalone_dma_fifo_wrport_we;
wire [128:0] main_genericstandalone_dma_fifo_wrport_dat_w;
wire main_genericstandalone_dma_fifo_do_read;
wire [6:0] main_genericstandalone_dma_fifo_rdport_adr;
wire [128:0] main_genericstandalone_dma_fifo_rdport_dat_r;
wire main_genericstandalone_dma_fifo_rdport_re;
wire [7:0] main_genericstandalone_dma_fifo_level1;
wire main_genericstandalone_dma_fifo_almost_empty;
wire [127:0] main_genericstandalone_dma_fifo_fifo_in_payload_data;
wire main_genericstandalone_dma_fifo_fifo_in_eop;
wire [127:0] main_genericstandalone_dma_fifo_fifo_out_payload_data;
wire main_genericstandalone_dma_fifo_fifo_out_eop;
reg main_genericstandalone_dma_fifo_recv_activated = 1'd0;
wire main_genericstandalone_dma_fifo_do_write;
wire main_genericstandalone_dma_rawslicer_sink_stb;
reg main_genericstandalone_dma_rawslicer_sink_ack;
wire main_genericstandalone_dma_rawslicer_sink_last;
wire main_genericstandalone_dma_rawslicer_sink_eop;
wire [127:0] main_genericstandalone_dma_rawslicer_sink_payload_data;
wire [615:0] main_genericstandalone_dma_rawslicer_source;
reg main_genericstandalone_dma_rawslicer_source_stb;
reg [6:0] main_genericstandalone_dma_rawslicer_source_consume;
reg main_genericstandalone_dma_rawslicer_flush;
reg main_genericstandalone_dma_rawslicer_flush_done;
reg [735:0] main_genericstandalone_dma_rawslicer_buf = 736'd0;
reg [6:0] main_genericstandalone_dma_rawslicer_level = 7'd0;
reg [6:0] main_genericstandalone_dma_rawslicer_next_level;
reg main_genericstandalone_dma_rawslicer_load_buf;
reg main_genericstandalone_dma_rawslicer_shift_buf;
reg main_genericstandalone_dma_reset = 1'd0;
reg main_genericstandalone_dma_record_converter_source_stb;
wire main_genericstandalone_dma_record_converter_source_ack;
reg main_genericstandalone_dma_record_converter_source_last = 1'd0;
reg main_genericstandalone_dma_record_converter_source_eop;
reg [7:0] main_genericstandalone_dma_record_converter_source_payload_length = 8'd0;
wire [23:0] main_genericstandalone_dma_record_converter_source_payload_channel;
wire [63:0] main_genericstandalone_dma_record_converter_source_payload_timestamp;
wire [7:0] main_genericstandalone_dma_record_converter_source_payload_address;
reg [511:0] main_genericstandalone_dma_record_converter_source_payload_data;
reg main_genericstandalone_dma_record_converter_end_marker_found;
reg main_genericstandalone_dma_record_converter_flush;
wire [7:0] main_genericstandalone_dma_record_converter_record_raw_length;
wire [23:0] main_genericstandalone_dma_record_converter_record_raw_channel;
wire [63:0] main_genericstandalone_dma_record_converter_record_raw_timestamp;
wire [7:0] main_genericstandalone_dma_record_converter_record_raw_address;
wire [511:0] main_genericstandalone_dma_record_converter_record_raw_data;
reg [63:0] main_genericstandalone_dma_time_offset_storage_full = 64'd0;
wire [63:0] main_genericstandalone_dma_time_offset_storage;
reg main_genericstandalone_dma_time_offset_re = 1'd0;
reg main_genericstandalone_dma_time_offset_source_stb = 1'd0;
wire main_genericstandalone_dma_time_offset_source_ack;
reg main_genericstandalone_dma_time_offset_source_last = 1'd0;
reg main_genericstandalone_dma_time_offset_source_eop = 1'd0;
reg [7:0] main_genericstandalone_dma_time_offset_source_payload_length = 8'd0;
reg [23:0] main_genericstandalone_dma_time_offset_source_payload_channel = 24'd0;
reg [63:0] main_genericstandalone_dma_time_offset_source_payload_timestamp = 64'd0;
reg [7:0] main_genericstandalone_dma_time_offset_source_payload_address = 8'd0;
reg [511:0] main_genericstandalone_dma_time_offset_source_payload_data = 512'd0;
wire main_genericstandalone_dma_time_offset_sink_stb;
wire main_genericstandalone_dma_time_offset_sink_ack;
wire main_genericstandalone_dma_time_offset_sink_last;
wire main_genericstandalone_dma_time_offset_sink_eop;
wire [7:0] main_genericstandalone_dma_time_offset_sink_payload_length;
wire [23:0] main_genericstandalone_dma_time_offset_sink_payload_channel;
wire [63:0] main_genericstandalone_dma_time_offset_sink_payload_timestamp;
wire [7:0] main_genericstandalone_dma_time_offset_sink_payload_address;
wire [511:0] main_genericstandalone_dma_time_offset_sink_payload_data;
wire main_genericstandalone_dma_cri_master_error_re;
wire [1:0] main_genericstandalone_dma_cri_master_error_r;
reg [1:0] main_genericstandalone_dma_cri_master_error_w = 2'd0;
reg [23:0] main_genericstandalone_dma_cri_master_error_channel_status = 24'd0;
reg [63:0] main_genericstandalone_dma_cri_master_error_timestamp_status = 64'd0;
reg [15:0] main_genericstandalone_dma_cri_master_error_address_status = 16'd0;
wire main_genericstandalone_dma_cri_master_sink_stb;
reg main_genericstandalone_dma_cri_master_sink_ack;
wire main_genericstandalone_dma_cri_master_sink_last;
wire main_genericstandalone_dma_cri_master_sink_eop;
wire [7:0] main_genericstandalone_dma_cri_master_sink_payload_length;
wire [23:0] main_genericstandalone_dma_cri_master_sink_payload_channel;
wire [63:0] main_genericstandalone_dma_cri_master_sink_payload_timestamp;
wire [7:0] main_genericstandalone_dma_cri_master_sink_payload_address;
wire [511:0] main_genericstandalone_dma_cri_master_sink_payload_data;
reg [1:0] main_genericstandalone_dma_cri_master_cri_cmd;
wire [23:0] main_genericstandalone_dma_cri_master_cri_chan_sel;
wire [63:0] main_genericstandalone_dma_cri_master_cri_o_timestamp;
wire [511:0] main_genericstandalone_dma_cri_master_cri_o_data;
wire [7:0] main_genericstandalone_dma_cri_master_cri_o_address;
wire [2:0] main_genericstandalone_dma_cri_master_cri_o_status;
wire main_genericstandalone_dma_cri_master_cri_o_buffer_space_valid;
wire [15:0] main_genericstandalone_dma_cri_master_cri_o_buffer_space;
reg [63:0] main_genericstandalone_dma_cri_master_cri_i_timeout = 64'd0;
wire [31:0] main_genericstandalone_dma_cri_master_cri_i_data;
wire [63:0] main_genericstandalone_dma_cri_master_cri_i_timestamp;
wire [3:0] main_genericstandalone_dma_cri_master_cri_i_status;
reg main_genericstandalone_dma_cri_master_busy;
reg main_genericstandalone_dma_cri_master_underflow_trigger;
reg main_genericstandalone_dma_cri_master_link_error_trigger;
wire [28:0] main_genericstandalone_interface0_csr_bus_adr;
wire [31:0] main_genericstandalone_interface0_csr_bus_dat_w;
reg [31:0] main_genericstandalone_interface0_csr_bus_dat_r = 32'd0;
wire [3:0] main_genericstandalone_interface0_csr_bus_sel;
wire main_genericstandalone_interface0_csr_bus_cyc;
wire main_genericstandalone_interface0_csr_bus_stb;
reg main_genericstandalone_interface0_csr_bus_ack = 1'd0;
wire main_genericstandalone_interface0_csr_bus_we;
wire [2:0] main_genericstandalone_interface0_csr_bus_cti;
wire [1:0] main_genericstandalone_interface0_csr_bus_bte;
reg main_genericstandalone_interface0_csr_bus_err = 1'd0;
wire main_genericstandalone_target0_re;
wire [31:0] main_genericstandalone_target0_r;
wire [31:0] main_genericstandalone_target0_w;
wire main_genericstandalone_o_data15_re;
wire [31:0] main_genericstandalone_o_data15_r;
wire [31:0] main_genericstandalone_o_data15_w;
wire main_genericstandalone_o_data14_re;
wire [31:0] main_genericstandalone_o_data14_r;
wire [31:0] main_genericstandalone_o_data14_w;
wire main_genericstandalone_o_data13_re;
wire [31:0] main_genericstandalone_o_data13_r;
wire [31:0] main_genericstandalone_o_data13_w;
wire main_genericstandalone_o_data12_re;
wire [31:0] main_genericstandalone_o_data12_r;
wire [31:0] main_genericstandalone_o_data12_w;
wire main_genericstandalone_o_data11_re;
wire [31:0] main_genericstandalone_o_data11_r;
wire [31:0] main_genericstandalone_o_data11_w;
wire main_genericstandalone_o_data10_re;
wire [31:0] main_genericstandalone_o_data10_r;
wire [31:0] main_genericstandalone_o_data10_w;
wire main_genericstandalone_o_data9_re;
wire [31:0] main_genericstandalone_o_data9_r;
wire [31:0] main_genericstandalone_o_data9_w;
wire main_genericstandalone_o_data8_re;
wire [31:0] main_genericstandalone_o_data8_r;
wire [31:0] main_genericstandalone_o_data8_w;
wire main_genericstandalone_o_data7_re;
wire [31:0] main_genericstandalone_o_data7_r;
wire [31:0] main_genericstandalone_o_data7_w;
wire main_genericstandalone_o_data6_re;
wire [31:0] main_genericstandalone_o_data6_r;
wire [31:0] main_genericstandalone_o_data6_w;
wire main_genericstandalone_o_data5_re;
wire [31:0] main_genericstandalone_o_data5_r;
wire [31:0] main_genericstandalone_o_data5_w;
wire main_genericstandalone_o_data4_re;
wire [31:0] main_genericstandalone_o_data4_r;
wire [31:0] main_genericstandalone_o_data4_w;
wire main_genericstandalone_o_data3_re;
wire [31:0] main_genericstandalone_o_data3_r;
wire [31:0] main_genericstandalone_o_data3_w;
wire main_genericstandalone_o_data2_re;
wire [31:0] main_genericstandalone_o_data2_r;
wire [31:0] main_genericstandalone_o_data2_w;
wire main_genericstandalone_o_data1_re;
wire [31:0] main_genericstandalone_o_data1_r;
wire [31:0] main_genericstandalone_o_data1_w;
wire main_genericstandalone_o_data0_re;
wire [31:0] main_genericstandalone_o_data0_r;
wire [31:0] main_genericstandalone_o_data0_w;
wire main_genericstandalone_o_status_re;
wire [2:0] main_genericstandalone_o_status_r;
wire [2:0] main_genericstandalone_o_status_w;
wire main_genericstandalone_i_timeout1_re;
wire [31:0] main_genericstandalone_i_timeout1_r;
wire [31:0] main_genericstandalone_i_timeout1_w;
wire main_genericstandalone_i_timeout0_re;
wire [31:0] main_genericstandalone_i_timeout0_r;
wire [31:0] main_genericstandalone_i_timeout0_w;
wire main_genericstandalone_i_data_re;
wire [31:0] main_genericstandalone_i_data_r;
wire [31:0] main_genericstandalone_i_data_w;
wire main_genericstandalone_i_timestamp1_re;
wire [31:0] main_genericstandalone_i_timestamp1_r;
wire [31:0] main_genericstandalone_i_timestamp1_w;
wire main_genericstandalone_i_timestamp0_re;
wire [31:0] main_genericstandalone_i_timestamp0_r;
wire [31:0] main_genericstandalone_i_timestamp0_w;
wire main_genericstandalone_i_status_re;
wire [3:0] main_genericstandalone_i_status_r;
wire [3:0] main_genericstandalone_i_status_w;
wire main_genericstandalone_counter1_re;
wire [31:0] main_genericstandalone_counter1_r;
wire [31:0] main_genericstandalone_counter1_w;
wire main_genericstandalone_counter0_re;
wire [31:0] main_genericstandalone_counter0_r;
wire [31:0] main_genericstandalone_counter0_w;
wire [28:0] main_genericstandalone_interface1_csr_bus_adr;
wire [31:0] main_genericstandalone_interface1_csr_bus_dat_w;
reg [31:0] main_genericstandalone_interface1_csr_bus_dat_r = 32'd0;
wire [3:0] main_genericstandalone_interface1_csr_bus_sel;
wire main_genericstandalone_interface1_csr_bus_cyc;
wire main_genericstandalone_interface1_csr_bus_stb;
reg main_genericstandalone_interface1_csr_bus_ack = 1'd0;
wire main_genericstandalone_interface1_csr_bus_we;
wire [2:0] main_genericstandalone_interface1_csr_bus_cti;
wire [1:0] main_genericstandalone_interface1_csr_bus_bte;
reg main_genericstandalone_interface1_csr_bus_err = 1'd0;
wire main_genericstandalone_base_address1_re;
wire main_genericstandalone_base_address1_r;
wire main_genericstandalone_base_address1_w;
wire main_genericstandalone_base_address0_re;
wire [31:0] main_genericstandalone_base_address0_r;
wire [31:0] main_genericstandalone_base_address0_w;
wire main_genericstandalone_time_offset1_re;
wire [31:0] main_genericstandalone_time_offset1_r;
wire [31:0] main_genericstandalone_time_offset1_w;
wire main_genericstandalone_time_offset0_re;
wire [31:0] main_genericstandalone_time_offset0_r;
wire [31:0] main_genericstandalone_time_offset0_w;
wire main_genericstandalone_error_channel_re;
wire [23:0] main_genericstandalone_error_channel_r;
wire [23:0] main_genericstandalone_error_channel_w;
wire main_genericstandalone_error_timestamp1_re;
wire [31:0] main_genericstandalone_error_timestamp1_r;
wire [31:0] main_genericstandalone_error_timestamp1_w;
wire main_genericstandalone_error_timestamp0_re;
wire [31:0] main_genericstandalone_error_timestamp0_r;
wire [31:0] main_genericstandalone_error_timestamp0_w;
wire main_genericstandalone_error_address_re;
wire [15:0] main_genericstandalone_error_address_r;
wire [15:0] main_genericstandalone_error_address_w;
wire [1:0] main_genericstandalone_cri_con_shared_cmd;
wire [23:0] main_genericstandalone_cri_con_shared_chan_sel;
wire [63:0] main_genericstandalone_cri_con_shared_o_timestamp;
wire [511:0] main_genericstandalone_cri_con_shared_o_data;
wire [7:0] main_genericstandalone_cri_con_shared_o_address;
reg [2:0] main_genericstandalone_cri_con_shared_o_status;
reg main_genericstandalone_cri_con_shared_o_buffer_space_valid;
reg [15:0] main_genericstandalone_cri_con_shared_o_buffer_space;
wire [63:0] main_genericstandalone_cri_con_shared_i_timeout;
reg [31:0] main_genericstandalone_cri_con_shared_i_data;
reg [63:0] main_genericstandalone_cri_con_shared_i_timestamp;
reg [3:0] main_genericstandalone_cri_con_shared_i_status;
reg [1:0] main_genericstandalone_cri_con_storage_full = 2'd0;
wire [1:0] main_genericstandalone_cri_con_storage;
reg main_genericstandalone_cri_con_re = 1'd0;
reg main_genericstandalone_cri_con_selected = 1'd0;
wire [28:0] main_genericstandalone_interface2_csr_bus_adr;
wire [31:0] main_genericstandalone_interface2_csr_bus_dat_w;
reg [31:0] main_genericstandalone_interface2_csr_bus_dat_r = 32'd0;
wire [3:0] main_genericstandalone_interface2_csr_bus_sel;
wire main_genericstandalone_interface2_csr_bus_cyc;
wire main_genericstandalone_interface2_csr_bus_stb;
reg main_genericstandalone_interface2_csr_bus_ack = 1'd0;
wire main_genericstandalone_interface2_csr_bus_we;
wire [2:0] main_genericstandalone_interface2_csr_bus_cti;
wire [1:0] main_genericstandalone_interface2_csr_bus_bte;
reg main_genericstandalone_interface2_csr_bus_err = 1'd0;
wire main_genericstandalone_selected0_re;
wire [1:0] main_genericstandalone_selected0_r;
wire [1:0] main_genericstandalone_selected0_w;
reg [5:0] main_genericstandalone_mon_chan_sel_storage_full = 6'd0;
wire [5:0] main_genericstandalone_mon_chan_sel_storage;
reg main_genericstandalone_mon_chan_sel_re = 1'd0;
reg [4:0] main_genericstandalone_mon_probe_sel_storage_full = 5'd0;
wire [4:0] main_genericstandalone_mon_probe_sel_storage;
reg main_genericstandalone_mon_probe_sel_re = 1'd0;
wire main_genericstandalone_mon_value_update_re;
wire main_genericstandalone_mon_value_update_r;
reg main_genericstandalone_mon_value_update_w = 1'd0;
reg [31:0] main_genericstandalone_mon_status = 32'd0;
wire main_genericstandalone_mon_bussynchronizer0_i;
wire main_genericstandalone_mon_bussynchronizer0_o;
wire main_genericstandalone_mon_bussynchronizer1_i;
wire main_genericstandalone_mon_bussynchronizer1_o;
wire main_genericstandalone_mon_bussynchronizer2_i;
wire main_genericstandalone_mon_bussynchronizer2_o;
wire main_genericstandalone_mon_bussynchronizer3_i;
wire main_genericstandalone_mon_bussynchronizer3_o;
wire main_genericstandalone_mon_bussynchronizer4_i;
wire main_genericstandalone_mon_bussynchronizer4_o;
wire main_genericstandalone_mon_bussynchronizer5_i;
wire main_genericstandalone_mon_bussynchronizer5_o;
wire main_genericstandalone_mon_bussynchronizer6_i;
wire main_genericstandalone_mon_bussynchronizer6_o;
wire main_genericstandalone_mon_bussynchronizer7_i;
wire main_genericstandalone_mon_bussynchronizer7_o;
wire main_genericstandalone_mon_bussynchronizer8_i;
wire main_genericstandalone_mon_bussynchronizer8_o;
wire main_genericstandalone_mon_bussynchronizer9_i;
wire main_genericstandalone_mon_bussynchronizer9_o;
wire main_genericstandalone_mon_bussynchronizer10_i;
wire main_genericstandalone_mon_bussynchronizer10_o;
wire main_genericstandalone_mon_bussynchronizer11_i;
wire main_genericstandalone_mon_bussynchronizer11_o;
wire main_genericstandalone_mon_bussynchronizer12_i;
wire main_genericstandalone_mon_bussynchronizer12_o;
wire main_genericstandalone_mon_bussynchronizer13_i;
wire main_genericstandalone_mon_bussynchronizer13_o;
wire main_genericstandalone_mon_bussynchronizer14_i;
wire main_genericstandalone_mon_bussynchronizer14_o;
wire main_genericstandalone_mon_bussynchronizer15_i;
wire main_genericstandalone_mon_bussynchronizer15_o;
wire main_genericstandalone_mon_bussynchronizer16_i;
wire main_genericstandalone_mon_bussynchronizer16_o;
wire main_genericstandalone_mon_bussynchronizer17_i;
wire main_genericstandalone_mon_bussynchronizer17_o;
wire main_genericstandalone_mon_bussynchronizer18_i;
wire main_genericstandalone_mon_bussynchronizer18_o;
wire main_genericstandalone_mon_bussynchronizer19_i;
wire main_genericstandalone_mon_bussynchronizer19_o;
wire [31:0] main_genericstandalone_mon_bussynchronizer20_i;
reg [31:0] main_genericstandalone_mon_bussynchronizer20_o = 32'd0;
reg main_genericstandalone_mon_bussynchronizer20_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer20_ping_i;
wire main_genericstandalone_mon_bussynchronizer20_ping_o0;
reg main_genericstandalone_mon_bussynchronizer20_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer20_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer20_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer20_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer20_pong_i;
wire main_genericstandalone_mon_bussynchronizer20_pong_o;
reg main_genericstandalone_mon_bussynchronizer20_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer20_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer20_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer20_wait;
wire main_genericstandalone_mon_bussynchronizer20_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer20_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_genericstandalone_mon_bussynchronizer20_ibuffer = 32'd0;
wire [31:0] main_genericstandalone_mon_bussynchronizer20_obuffer;
wire [31:0] main_genericstandalone_mon_bussynchronizer21_i;
reg [31:0] main_genericstandalone_mon_bussynchronizer21_o = 32'd0;
reg main_genericstandalone_mon_bussynchronizer21_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer21_ping_i;
wire main_genericstandalone_mon_bussynchronizer21_ping_o0;
reg main_genericstandalone_mon_bussynchronizer21_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer21_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer21_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer21_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer21_pong_i;
wire main_genericstandalone_mon_bussynchronizer21_pong_o;
reg main_genericstandalone_mon_bussynchronizer21_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer21_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer21_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer21_wait;
wire main_genericstandalone_mon_bussynchronizer21_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer21_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_genericstandalone_mon_bussynchronizer21_ibuffer = 32'd0;
wire [31:0] main_genericstandalone_mon_bussynchronizer21_obuffer;
wire [31:0] main_genericstandalone_mon_bussynchronizer22_i;
reg [31:0] main_genericstandalone_mon_bussynchronizer22_o = 32'd0;
reg main_genericstandalone_mon_bussynchronizer22_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer22_ping_i;
wire main_genericstandalone_mon_bussynchronizer22_ping_o0;
reg main_genericstandalone_mon_bussynchronizer22_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer22_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer22_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer22_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer22_pong_i;
wire main_genericstandalone_mon_bussynchronizer22_pong_o;
reg main_genericstandalone_mon_bussynchronizer22_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer22_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer22_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer22_wait;
wire main_genericstandalone_mon_bussynchronizer22_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer22_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_genericstandalone_mon_bussynchronizer22_ibuffer = 32'd0;
wire [31:0] main_genericstandalone_mon_bussynchronizer22_obuffer;
wire [31:0] main_genericstandalone_mon_bussynchronizer23_i;
reg [31:0] main_genericstandalone_mon_bussynchronizer23_o = 32'd0;
reg main_genericstandalone_mon_bussynchronizer23_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer23_ping_i;
wire main_genericstandalone_mon_bussynchronizer23_ping_o0;
reg main_genericstandalone_mon_bussynchronizer23_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer23_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer23_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer23_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer23_pong_i;
wire main_genericstandalone_mon_bussynchronizer23_pong_o;
reg main_genericstandalone_mon_bussynchronizer23_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer23_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer23_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer23_wait;
wire main_genericstandalone_mon_bussynchronizer23_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer23_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_genericstandalone_mon_bussynchronizer23_ibuffer = 32'd0;
wire [31:0] main_genericstandalone_mon_bussynchronizer23_obuffer;
wire main_genericstandalone_mon_bussynchronizer24_i;
wire main_genericstandalone_mon_bussynchronizer24_o;
wire main_genericstandalone_mon_bussynchronizer25_i;
wire main_genericstandalone_mon_bussynchronizer25_o;
wire main_genericstandalone_mon_bussynchronizer26_i;
wire main_genericstandalone_mon_bussynchronizer26_o;
wire main_genericstandalone_mon_bussynchronizer27_i;
wire main_genericstandalone_mon_bussynchronizer27_o;
wire main_genericstandalone_mon_bussynchronizer28_i;
wire main_genericstandalone_mon_bussynchronizer28_o;
wire [31:0] main_genericstandalone_mon_bussynchronizer29_i;
reg [31:0] main_genericstandalone_mon_bussynchronizer29_o = 32'd0;
reg main_genericstandalone_mon_bussynchronizer29_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer29_ping_i;
wire main_genericstandalone_mon_bussynchronizer29_ping_o0;
reg main_genericstandalone_mon_bussynchronizer29_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer29_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer29_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer29_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer29_pong_i;
wire main_genericstandalone_mon_bussynchronizer29_pong_o;
reg main_genericstandalone_mon_bussynchronizer29_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer29_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer29_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer29_wait;
wire main_genericstandalone_mon_bussynchronizer29_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer29_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_genericstandalone_mon_bussynchronizer29_ibuffer = 32'd0;
wire [31:0] main_genericstandalone_mon_bussynchronizer29_obuffer;
wire [31:0] main_genericstandalone_mon_bussynchronizer30_i;
reg [31:0] main_genericstandalone_mon_bussynchronizer30_o = 32'd0;
reg main_genericstandalone_mon_bussynchronizer30_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer30_ping_i;
wire main_genericstandalone_mon_bussynchronizer30_ping_o0;
reg main_genericstandalone_mon_bussynchronizer30_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer30_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer30_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer30_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer30_pong_i;
wire main_genericstandalone_mon_bussynchronizer30_pong_o;
reg main_genericstandalone_mon_bussynchronizer30_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer30_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer30_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer30_wait;
wire main_genericstandalone_mon_bussynchronizer30_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer30_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_genericstandalone_mon_bussynchronizer30_ibuffer = 32'd0;
wire [31:0] main_genericstandalone_mon_bussynchronizer30_obuffer;
wire [31:0] main_genericstandalone_mon_bussynchronizer31_i;
reg [31:0] main_genericstandalone_mon_bussynchronizer31_o = 32'd0;
reg main_genericstandalone_mon_bussynchronizer31_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer31_ping_i;
wire main_genericstandalone_mon_bussynchronizer31_ping_o0;
reg main_genericstandalone_mon_bussynchronizer31_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer31_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer31_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer31_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer31_pong_i;
wire main_genericstandalone_mon_bussynchronizer31_pong_o;
reg main_genericstandalone_mon_bussynchronizer31_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer31_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer31_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer31_wait;
wire main_genericstandalone_mon_bussynchronizer31_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer31_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_genericstandalone_mon_bussynchronizer31_ibuffer = 32'd0;
wire [31:0] main_genericstandalone_mon_bussynchronizer31_obuffer;
wire [31:0] main_genericstandalone_mon_bussynchronizer32_i;
reg [31:0] main_genericstandalone_mon_bussynchronizer32_o = 32'd0;
reg main_genericstandalone_mon_bussynchronizer32_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer32_ping_i;
wire main_genericstandalone_mon_bussynchronizer32_ping_o0;
reg main_genericstandalone_mon_bussynchronizer32_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer32_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer32_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer32_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer32_pong_i;
wire main_genericstandalone_mon_bussynchronizer32_pong_o;
reg main_genericstandalone_mon_bussynchronizer32_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer32_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer32_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer32_wait;
wire main_genericstandalone_mon_bussynchronizer32_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer32_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_genericstandalone_mon_bussynchronizer32_ibuffer = 32'd0;
wire [31:0] main_genericstandalone_mon_bussynchronizer32_obuffer;
wire main_genericstandalone_mon_bussynchronizer33_i;
wire main_genericstandalone_mon_bussynchronizer33_o;
wire main_genericstandalone_mon_bussynchronizer34_i;
wire main_genericstandalone_mon_bussynchronizer34_o;
wire main_genericstandalone_mon_bussynchronizer35_i;
wire main_genericstandalone_mon_bussynchronizer35_o;
wire main_genericstandalone_mon_bussynchronizer36_i;
wire main_genericstandalone_mon_bussynchronizer36_o;
wire main_genericstandalone_mon_bussynchronizer37_i;
wire main_genericstandalone_mon_bussynchronizer37_o;
wire main_genericstandalone_mon_bussynchronizer38_i;
wire main_genericstandalone_mon_bussynchronizer38_o;
wire [15:0] main_genericstandalone_mon_bussynchronizer39_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer39_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer39_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer39_ping_i;
wire main_genericstandalone_mon_bussynchronizer39_ping_o0;
reg main_genericstandalone_mon_bussynchronizer39_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer39_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer39_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer39_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer39_pong_i;
wire main_genericstandalone_mon_bussynchronizer39_pong_o;
reg main_genericstandalone_mon_bussynchronizer39_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer39_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer39_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer39_wait;
wire main_genericstandalone_mon_bussynchronizer39_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer39_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer39_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer39_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer40_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer40_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer40_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer40_ping_i;
wire main_genericstandalone_mon_bussynchronizer40_ping_o0;
reg main_genericstandalone_mon_bussynchronizer40_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer40_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer40_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer40_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer40_pong_i;
wire main_genericstandalone_mon_bussynchronizer40_pong_o;
reg main_genericstandalone_mon_bussynchronizer40_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer40_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer40_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer40_wait;
wire main_genericstandalone_mon_bussynchronizer40_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer40_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer40_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer40_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer41_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer41_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer41_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer41_ping_i;
wire main_genericstandalone_mon_bussynchronizer41_ping_o0;
reg main_genericstandalone_mon_bussynchronizer41_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer41_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer41_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer41_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer41_pong_i;
wire main_genericstandalone_mon_bussynchronizer41_pong_o;
reg main_genericstandalone_mon_bussynchronizer41_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer41_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer41_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer41_wait;
wire main_genericstandalone_mon_bussynchronizer41_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer41_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer41_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer41_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer42_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer42_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer42_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer42_ping_i;
wire main_genericstandalone_mon_bussynchronizer42_ping_o0;
reg main_genericstandalone_mon_bussynchronizer42_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer42_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer42_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer42_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer42_pong_i;
wire main_genericstandalone_mon_bussynchronizer42_pong_o;
reg main_genericstandalone_mon_bussynchronizer42_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer42_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer42_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer42_wait;
wire main_genericstandalone_mon_bussynchronizer42_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer42_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer42_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer42_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer43_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer43_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer43_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer43_ping_i;
wire main_genericstandalone_mon_bussynchronizer43_ping_o0;
reg main_genericstandalone_mon_bussynchronizer43_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer43_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer43_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer43_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer43_pong_i;
wire main_genericstandalone_mon_bussynchronizer43_pong_o;
reg main_genericstandalone_mon_bussynchronizer43_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer43_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer43_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer43_wait;
wire main_genericstandalone_mon_bussynchronizer43_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer43_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer43_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer43_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer44_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer44_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer44_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer44_ping_i;
wire main_genericstandalone_mon_bussynchronizer44_ping_o0;
reg main_genericstandalone_mon_bussynchronizer44_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer44_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer44_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer44_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer44_pong_i;
wire main_genericstandalone_mon_bussynchronizer44_pong_o;
reg main_genericstandalone_mon_bussynchronizer44_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer44_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer44_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer44_wait;
wire main_genericstandalone_mon_bussynchronizer44_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer44_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer44_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer44_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer45_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer45_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer45_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer45_ping_i;
wire main_genericstandalone_mon_bussynchronizer45_ping_o0;
reg main_genericstandalone_mon_bussynchronizer45_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer45_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer45_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer45_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer45_pong_i;
wire main_genericstandalone_mon_bussynchronizer45_pong_o;
reg main_genericstandalone_mon_bussynchronizer45_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer45_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer45_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer45_wait;
wire main_genericstandalone_mon_bussynchronizer45_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer45_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer45_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer45_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer46_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer46_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer46_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer46_ping_i;
wire main_genericstandalone_mon_bussynchronizer46_ping_o0;
reg main_genericstandalone_mon_bussynchronizer46_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer46_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer46_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer46_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer46_pong_i;
wire main_genericstandalone_mon_bussynchronizer46_pong_o;
reg main_genericstandalone_mon_bussynchronizer46_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer46_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer46_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer46_wait;
wire main_genericstandalone_mon_bussynchronizer46_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer46_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer46_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer46_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer47_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer47_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer47_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer47_ping_i;
wire main_genericstandalone_mon_bussynchronizer47_ping_o0;
reg main_genericstandalone_mon_bussynchronizer47_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer47_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer47_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer47_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer47_pong_i;
wire main_genericstandalone_mon_bussynchronizer47_pong_o;
reg main_genericstandalone_mon_bussynchronizer47_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer47_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer47_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer47_wait;
wire main_genericstandalone_mon_bussynchronizer47_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer47_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer47_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer47_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer48_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer48_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer48_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer48_ping_i;
wire main_genericstandalone_mon_bussynchronizer48_ping_o0;
reg main_genericstandalone_mon_bussynchronizer48_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer48_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer48_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer48_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer48_pong_i;
wire main_genericstandalone_mon_bussynchronizer48_pong_o;
reg main_genericstandalone_mon_bussynchronizer48_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer48_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer48_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer48_wait;
wire main_genericstandalone_mon_bussynchronizer48_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer48_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer48_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer48_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer49_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer49_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer49_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer49_ping_i;
wire main_genericstandalone_mon_bussynchronizer49_ping_o0;
reg main_genericstandalone_mon_bussynchronizer49_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer49_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer49_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer49_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer49_pong_i;
wire main_genericstandalone_mon_bussynchronizer49_pong_o;
reg main_genericstandalone_mon_bussynchronizer49_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer49_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer49_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer49_wait;
wire main_genericstandalone_mon_bussynchronizer49_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer49_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer49_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer49_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer50_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer50_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer50_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer50_ping_i;
wire main_genericstandalone_mon_bussynchronizer50_ping_o0;
reg main_genericstandalone_mon_bussynchronizer50_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer50_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer50_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer50_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer50_pong_i;
wire main_genericstandalone_mon_bussynchronizer50_pong_o;
reg main_genericstandalone_mon_bussynchronizer50_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer50_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer50_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer50_wait;
wire main_genericstandalone_mon_bussynchronizer50_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer50_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer50_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer50_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer51_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer51_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer51_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer51_ping_i;
wire main_genericstandalone_mon_bussynchronizer51_ping_o0;
reg main_genericstandalone_mon_bussynchronizer51_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer51_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer51_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer51_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer51_pong_i;
wire main_genericstandalone_mon_bussynchronizer51_pong_o;
reg main_genericstandalone_mon_bussynchronizer51_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer51_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer51_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer51_wait;
wire main_genericstandalone_mon_bussynchronizer51_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer51_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer51_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer51_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer52_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer52_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer52_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer52_ping_i;
wire main_genericstandalone_mon_bussynchronizer52_ping_o0;
reg main_genericstandalone_mon_bussynchronizer52_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer52_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer52_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer52_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer52_pong_i;
wire main_genericstandalone_mon_bussynchronizer52_pong_o;
reg main_genericstandalone_mon_bussynchronizer52_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer52_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer52_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer52_wait;
wire main_genericstandalone_mon_bussynchronizer52_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer52_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer52_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer52_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer53_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer53_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer53_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer53_ping_i;
wire main_genericstandalone_mon_bussynchronizer53_ping_o0;
reg main_genericstandalone_mon_bussynchronizer53_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer53_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer53_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer53_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer53_pong_i;
wire main_genericstandalone_mon_bussynchronizer53_pong_o;
reg main_genericstandalone_mon_bussynchronizer53_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer53_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer53_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer53_wait;
wire main_genericstandalone_mon_bussynchronizer53_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer53_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer53_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer53_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer54_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer54_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer54_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer54_ping_i;
wire main_genericstandalone_mon_bussynchronizer54_ping_o0;
reg main_genericstandalone_mon_bussynchronizer54_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer54_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer54_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer54_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer54_pong_i;
wire main_genericstandalone_mon_bussynchronizer54_pong_o;
reg main_genericstandalone_mon_bussynchronizer54_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer54_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer54_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer54_wait;
wire main_genericstandalone_mon_bussynchronizer54_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer54_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer54_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer54_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer55_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer55_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer55_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer55_ping_i;
wire main_genericstandalone_mon_bussynchronizer55_ping_o0;
reg main_genericstandalone_mon_bussynchronizer55_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer55_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer55_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer55_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer55_pong_i;
wire main_genericstandalone_mon_bussynchronizer55_pong_o;
reg main_genericstandalone_mon_bussynchronizer55_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer55_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer55_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer55_wait;
wire main_genericstandalone_mon_bussynchronizer55_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer55_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer55_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer55_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer56_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer56_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer56_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer56_ping_i;
wire main_genericstandalone_mon_bussynchronizer56_ping_o0;
reg main_genericstandalone_mon_bussynchronizer56_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer56_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer56_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer56_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer56_pong_i;
wire main_genericstandalone_mon_bussynchronizer56_pong_o;
reg main_genericstandalone_mon_bussynchronizer56_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer56_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer56_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer56_wait;
wire main_genericstandalone_mon_bussynchronizer56_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer56_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer56_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer56_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer57_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer57_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer57_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer57_ping_i;
wire main_genericstandalone_mon_bussynchronizer57_ping_o0;
reg main_genericstandalone_mon_bussynchronizer57_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer57_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer57_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer57_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer57_pong_i;
wire main_genericstandalone_mon_bussynchronizer57_pong_o;
reg main_genericstandalone_mon_bussynchronizer57_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer57_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer57_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer57_wait;
wire main_genericstandalone_mon_bussynchronizer57_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer57_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer57_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer57_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer58_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer58_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer58_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer58_ping_i;
wire main_genericstandalone_mon_bussynchronizer58_ping_o0;
reg main_genericstandalone_mon_bussynchronizer58_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer58_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer58_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer58_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer58_pong_i;
wire main_genericstandalone_mon_bussynchronizer58_pong_o;
reg main_genericstandalone_mon_bussynchronizer58_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer58_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer58_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer58_wait;
wire main_genericstandalone_mon_bussynchronizer58_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer58_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer58_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer58_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer59_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer59_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer59_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer59_ping_i;
wire main_genericstandalone_mon_bussynchronizer59_ping_o0;
reg main_genericstandalone_mon_bussynchronizer59_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer59_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer59_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer59_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer59_pong_i;
wire main_genericstandalone_mon_bussynchronizer59_pong_o;
reg main_genericstandalone_mon_bussynchronizer59_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer59_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer59_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer59_wait;
wire main_genericstandalone_mon_bussynchronizer59_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer59_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer59_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer59_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer60_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer60_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer60_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer60_ping_i;
wire main_genericstandalone_mon_bussynchronizer60_ping_o0;
reg main_genericstandalone_mon_bussynchronizer60_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer60_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer60_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer60_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer60_pong_i;
wire main_genericstandalone_mon_bussynchronizer60_pong_o;
reg main_genericstandalone_mon_bussynchronizer60_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer60_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer60_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer60_wait;
wire main_genericstandalone_mon_bussynchronizer60_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer60_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer60_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer60_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer61_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer61_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer61_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer61_ping_i;
wire main_genericstandalone_mon_bussynchronizer61_ping_o0;
reg main_genericstandalone_mon_bussynchronizer61_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer61_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer61_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer61_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer61_pong_i;
wire main_genericstandalone_mon_bussynchronizer61_pong_o;
reg main_genericstandalone_mon_bussynchronizer61_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer61_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer61_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer61_wait;
wire main_genericstandalone_mon_bussynchronizer61_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer61_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer61_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer61_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer62_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer62_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer62_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer62_ping_i;
wire main_genericstandalone_mon_bussynchronizer62_ping_o0;
reg main_genericstandalone_mon_bussynchronizer62_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer62_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer62_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer62_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer62_pong_i;
wire main_genericstandalone_mon_bussynchronizer62_pong_o;
reg main_genericstandalone_mon_bussynchronizer62_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer62_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer62_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer62_wait;
wire main_genericstandalone_mon_bussynchronizer62_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer62_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer62_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer62_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer63_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer63_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer63_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer63_ping_i;
wire main_genericstandalone_mon_bussynchronizer63_ping_o0;
reg main_genericstandalone_mon_bussynchronizer63_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer63_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer63_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer63_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer63_pong_i;
wire main_genericstandalone_mon_bussynchronizer63_pong_o;
reg main_genericstandalone_mon_bussynchronizer63_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer63_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer63_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer63_wait;
wire main_genericstandalone_mon_bussynchronizer63_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer63_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer63_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer63_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer64_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer64_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer64_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer64_ping_i;
wire main_genericstandalone_mon_bussynchronizer64_ping_o0;
reg main_genericstandalone_mon_bussynchronizer64_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer64_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer64_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer64_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer64_pong_i;
wire main_genericstandalone_mon_bussynchronizer64_pong_o;
reg main_genericstandalone_mon_bussynchronizer64_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer64_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer64_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer64_wait;
wire main_genericstandalone_mon_bussynchronizer64_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer64_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer64_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer64_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer65_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer65_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer65_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer65_ping_i;
wire main_genericstandalone_mon_bussynchronizer65_ping_o0;
reg main_genericstandalone_mon_bussynchronizer65_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer65_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer65_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer65_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer65_pong_i;
wire main_genericstandalone_mon_bussynchronizer65_pong_o;
reg main_genericstandalone_mon_bussynchronizer65_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer65_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer65_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer65_wait;
wire main_genericstandalone_mon_bussynchronizer65_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer65_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer65_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer65_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer66_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer66_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer66_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer66_ping_i;
wire main_genericstandalone_mon_bussynchronizer66_ping_o0;
reg main_genericstandalone_mon_bussynchronizer66_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer66_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer66_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer66_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer66_pong_i;
wire main_genericstandalone_mon_bussynchronizer66_pong_o;
reg main_genericstandalone_mon_bussynchronizer66_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer66_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer66_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer66_wait;
wire main_genericstandalone_mon_bussynchronizer66_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer66_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer66_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer66_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer67_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer67_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer67_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer67_ping_i;
wire main_genericstandalone_mon_bussynchronizer67_ping_o0;
reg main_genericstandalone_mon_bussynchronizer67_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer67_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer67_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer67_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer67_pong_i;
wire main_genericstandalone_mon_bussynchronizer67_pong_o;
reg main_genericstandalone_mon_bussynchronizer67_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer67_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer67_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer67_wait;
wire main_genericstandalone_mon_bussynchronizer67_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer67_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer67_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer67_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer68_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer68_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer68_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer68_ping_i;
wire main_genericstandalone_mon_bussynchronizer68_ping_o0;
reg main_genericstandalone_mon_bussynchronizer68_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer68_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer68_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer68_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer68_pong_i;
wire main_genericstandalone_mon_bussynchronizer68_pong_o;
reg main_genericstandalone_mon_bussynchronizer68_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer68_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer68_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer68_wait;
wire main_genericstandalone_mon_bussynchronizer68_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer68_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer68_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer68_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer69_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer69_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer69_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer69_ping_i;
wire main_genericstandalone_mon_bussynchronizer69_ping_o0;
reg main_genericstandalone_mon_bussynchronizer69_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer69_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer69_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer69_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer69_pong_i;
wire main_genericstandalone_mon_bussynchronizer69_pong_o;
reg main_genericstandalone_mon_bussynchronizer69_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer69_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer69_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer69_wait;
wire main_genericstandalone_mon_bussynchronizer69_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer69_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer69_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer69_obuffer;
wire [15:0] main_genericstandalone_mon_bussynchronizer70_i;
reg [15:0] main_genericstandalone_mon_bussynchronizer70_o = 16'd0;
reg main_genericstandalone_mon_bussynchronizer70_starter = 1'd1;
wire main_genericstandalone_mon_bussynchronizer70_ping_i;
wire main_genericstandalone_mon_bussynchronizer70_ping_o0;
reg main_genericstandalone_mon_bussynchronizer70_ping_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer70_ping_toggle_o;
reg main_genericstandalone_mon_bussynchronizer70_ping_toggle_o_r = 1'd0;
reg main_genericstandalone_mon_bussynchronizer70_ping_o1 = 1'd0;
wire main_genericstandalone_mon_bussynchronizer70_pong_i;
wire main_genericstandalone_mon_bussynchronizer70_pong_o;
reg main_genericstandalone_mon_bussynchronizer70_pong_toggle_i = 1'd0;
wire main_genericstandalone_mon_bussynchronizer70_pong_toggle_o;
reg main_genericstandalone_mon_bussynchronizer70_pong_toggle_o_r = 1'd0;
wire main_genericstandalone_mon_bussynchronizer70_wait;
wire main_genericstandalone_mon_bussynchronizer70_done;
reg [7:0] main_genericstandalone_mon_bussynchronizer70_count = 8'd128;
(* dont_touch = "true" *) reg [15:0] main_genericstandalone_mon_bussynchronizer70_ibuffer = 16'd0;
wire [15:0] main_genericstandalone_mon_bussynchronizer70_obuffer;
wire main_genericstandalone_mon_bussynchronizer71_i;
wire main_genericstandalone_mon_bussynchronizer71_o;
wire main_genericstandalone_mon_bussynchronizer72_i;
wire main_genericstandalone_mon_bussynchronizer72_o;
wire main_genericstandalone_mon_bussynchronizer73_i;
wire main_genericstandalone_mon_bussynchronizer73_o;
wire main_genericstandalone_mon_bussynchronizer74_i;
wire main_genericstandalone_mon_bussynchronizer74_o;
wire main_genericstandalone_mon_bussynchronizer75_i;
wire main_genericstandalone_mon_bussynchronizer75_o;
reg [5:0] main_genericstandalone_inj_chan_sel_storage_full = 6'd0;
wire [5:0] main_genericstandalone_inj_chan_sel_storage;
reg main_genericstandalone_inj_chan_sel_re = 1'd0;
reg [1:0] main_genericstandalone_inj_override_sel_storage_full = 2'd0;
wire [1:0] main_genericstandalone_inj_override_sel_storage;
reg main_genericstandalone_inj_override_sel_re = 1'd0;
wire main_genericstandalone_inj_value_re;
wire main_genericstandalone_inj_value_r;
wire main_genericstandalone_inj_value_w;
reg main_genericstandalone_inj_o_sys0 = 1'd0;
reg main_genericstandalone_inj_o_sys1 = 1'd0;
reg main_genericstandalone_inj_o_sys2 = 1'd0;
reg main_genericstandalone_inj_o_sys3 = 1'd0;
reg main_genericstandalone_inj_o_sys4 = 1'd0;
reg main_genericstandalone_inj_o_sys5 = 1'd0;
reg main_genericstandalone_inj_o_sys6 = 1'd0;
reg main_genericstandalone_inj_o_sys7 = 1'd0;
reg main_genericstandalone_inj_o_sys8 = 1'd0;
reg main_genericstandalone_inj_o_sys9 = 1'd0;
reg main_genericstandalone_inj_o_sys10 = 1'd0;
reg main_genericstandalone_inj_o_sys11 = 1'd0;
reg main_genericstandalone_inj_o_sys12 = 1'd0;
reg main_genericstandalone_inj_o_sys13 = 1'd0;
reg main_genericstandalone_inj_o_sys14 = 1'd0;
reg main_genericstandalone_inj_o_sys15 = 1'd0;
reg main_genericstandalone_inj_o_sys16 = 1'd0;
reg main_genericstandalone_inj_o_sys17 = 1'd0;
reg main_genericstandalone_inj_o_sys18 = 1'd0;
reg main_genericstandalone_inj_o_sys19 = 1'd0;
reg main_genericstandalone_inj_o_sys20 = 1'd0;
reg main_genericstandalone_inj_o_sys21 = 1'd0;
reg main_genericstandalone_inj_o_sys22 = 1'd0;
reg main_genericstandalone_inj_o_sys23 = 1'd0;
reg main_genericstandalone_inj_o_sys24 = 1'd0;
reg main_genericstandalone_inj_o_sys25 = 1'd0;
reg main_genericstandalone_inj_o_sys26 = 1'd0;
reg main_genericstandalone_inj_o_sys27 = 1'd0;
reg main_genericstandalone_inj_o_sys28 = 1'd0;
reg main_genericstandalone_inj_o_sys29 = 1'd0;
reg main_genericstandalone_inj_o_sys30 = 1'd0;
reg main_genericstandalone_inj_o_sys31 = 1'd0;
reg main_genericstandalone_inj_o_sys32 = 1'd0;
reg main_genericstandalone_inj_o_sys33 = 1'd0;
reg main_genericstandalone_inj_o_sys34 = 1'd0;
reg main_genericstandalone_inj_o_sys35 = 1'd0;
reg main_genericstandalone_inj_o_sys36 = 1'd0;
reg main_genericstandalone_inj_o_sys37 = 1'd0;
reg main_genericstandalone_inj_o_sys38 = 1'd0;
reg main_genericstandalone_inj_o_sys39 = 1'd0;
reg main_genericstandalone_inj_o_sys40 = 1'd0;
reg main_genericstandalone_inj_o_sys41 = 1'd0;
reg main_genericstandalone_inj_o_sys42 = 1'd0;
reg main_genericstandalone_inj_o_sys43 = 1'd0;
reg main_genericstandalone_inj_o_sys44 = 1'd0;
reg main_genericstandalone_inj_o_sys45 = 1'd0;
reg main_genericstandalone_inj_o_sys46 = 1'd0;
reg main_genericstandalone_inj_o_sys47 = 1'd0;
reg main_genericstandalone_inj_o_sys48 = 1'd0;
reg main_genericstandalone_inj_o_sys49 = 1'd0;
reg main_genericstandalone_inj_o_sys50 = 1'd0;
reg main_genericstandalone_inj_o_sys51 = 1'd0;
reg main_genericstandalone_inj_o_sys52 = 1'd0;
reg main_genericstandalone_inj_o_sys53 = 1'd0;
reg main_genericstandalone_inj_o_sys54 = 1'd0;
reg main_genericstandalone_inj_o_sys55 = 1'd0;
reg main_genericstandalone_inj_o_sys56 = 1'd0;
reg main_genericstandalone_inj_o_sys57 = 1'd0;
reg main_genericstandalone_inj_o_sys58 = 1'd0;
reg main_genericstandalone_inj_o_sys59 = 1'd0;
reg main_genericstandalone_inj_o_sys60 = 1'd0;
reg main_genericstandalone_inj_o_sys61 = 1'd0;
reg main_genericstandalone_inj_o_sys62 = 1'd0;
reg main_genericstandalone_inj_o_sys63 = 1'd0;
reg main_genericstandalone_inj_o_sys64 = 1'd0;
reg main_genericstandalone_inj_o_sys65 = 1'd0;
reg main_genericstandalone_inj_o_sys66 = 1'd0;
reg main_genericstandalone_inj_o_sys67 = 1'd0;
reg [28:0] main_genericstandalone_interface1_bus_adr = 29'd0;
wire [127:0] main_genericstandalone_interface1_bus_dat_w;
wire [127:0] main_genericstandalone_interface1_bus_dat_r;
wire [15:0] main_genericstandalone_interface1_bus_sel;
wire main_genericstandalone_interface1_bus_cyc;
wire main_genericstandalone_interface1_bus_stb;
wire main_genericstandalone_interface1_bus_ack;
wire main_genericstandalone_interface1_bus_we;
wire [2:0] main_genericstandalone_interface1_bus_cti;
reg [1:0] main_genericstandalone_interface1_bus_bte = 2'd0;
wire main_genericstandalone_interface1_bus_err;
reg main_genericstandalone_rtio_analyzer_enable_storage_full = 1'd0;
wire main_genericstandalone_rtio_analyzer_enable_storage;
reg main_genericstandalone_rtio_analyzer_enable_re = 1'd0;
reg main_genericstandalone_rtio_analyzer_busy_status = 1'd0;
reg main_genericstandalone_rtio_analyzer_message_encoder_source_stb = 1'd0;
wire main_genericstandalone_rtio_analyzer_message_encoder_source_ack;
reg main_genericstandalone_rtio_analyzer_message_encoder_source_last = 1'd0;
reg main_genericstandalone_rtio_analyzer_message_encoder_source_eop = 1'd0;
reg [255:0] main_genericstandalone_rtio_analyzer_message_encoder_source_payload_data = 256'd0;
reg main_genericstandalone_rtio_analyzer_message_encoder_status = 1'd0;
wire main_genericstandalone_rtio_analyzer_message_encoder_overflow_reset_re;
wire main_genericstandalone_rtio_analyzer_message_encoder_overflow_reset_r;
reg main_genericstandalone_rtio_analyzer_message_encoder_overflow_reset_w = 1'd0;
reg main_genericstandalone_rtio_analyzer_message_encoder_read_wait_event_r = 1'd0;
reg main_genericstandalone_rtio_analyzer_message_encoder_read_done;
reg main_genericstandalone_rtio_analyzer_message_encoder_read_overflow;
wire main_genericstandalone_rtio_analyzer_message_encoder_input_output_stb;
reg [1:0] main_genericstandalone_rtio_analyzer_message_encoder_input_output_message_type;
wire [29:0] main_genericstandalone_rtio_analyzer_message_encoder_input_output_channel;
reg [63:0] main_genericstandalone_rtio_analyzer_message_encoder_input_output_timestamp;
wire [63:0] main_genericstandalone_rtio_analyzer_message_encoder_input_output_rtio_counter;
wire [31:0] main_genericstandalone_rtio_analyzer_message_encoder_input_output_address_padding;
reg [63:0] main_genericstandalone_rtio_analyzer_message_encoder_input_output_data;
reg main_genericstandalone_rtio_analyzer_message_encoder_exception_stb;
wire [1:0] main_genericstandalone_rtio_analyzer_message_encoder_exception_message_type;
wire [29:0] main_genericstandalone_rtio_analyzer_message_encoder_exception_channel;
reg [63:0] main_genericstandalone_rtio_analyzer_message_encoder_exception_padding0 = 64'd0;
wire [63:0] main_genericstandalone_rtio_analyzer_message_encoder_exception_rtio_counter;
reg [7:0] main_genericstandalone_rtio_analyzer_message_encoder_exception_exception_type;
reg [87:0] main_genericstandalone_rtio_analyzer_message_encoder_exception_padding1 = 88'd0;
reg main_genericstandalone_rtio_analyzer_message_encoder_just_written = 1'd0;
wire [1:0] main_genericstandalone_rtio_analyzer_message_encoder_stopped_message_type;
reg [93:0] main_genericstandalone_rtio_analyzer_message_encoder_stopped_padding0 = 94'd0;
wire [63:0] main_genericstandalone_rtio_analyzer_message_encoder_stopped_rtio_counter;
reg [95:0] main_genericstandalone_rtio_analyzer_message_encoder_stopped_padding1 = 96'd0;
reg main_genericstandalone_rtio_analyzer_message_encoder_enable_r = 1'd0;
reg main_genericstandalone_rtio_analyzer_message_encoder_stopping = 1'd0;
wire main_genericstandalone_rtio_analyzer_fifo_sink_stb;
wire main_genericstandalone_rtio_analyzer_fifo_sink_ack;
wire main_genericstandalone_rtio_analyzer_fifo_sink_last;
wire main_genericstandalone_rtio_analyzer_fifo_sink_eop;
wire [255:0] main_genericstandalone_rtio_analyzer_fifo_sink_payload_data;
reg main_genericstandalone_rtio_analyzer_fifo_source_stb;
wire main_genericstandalone_rtio_analyzer_fifo_source_ack;
wire main_genericstandalone_rtio_analyzer_fifo_source_last;
wire main_genericstandalone_rtio_analyzer_fifo_source_eop;
wire [255:0] main_genericstandalone_rtio_analyzer_fifo_source_payload_data;
reg main_genericstandalone_rtio_analyzer_fifo_re;
reg main_genericstandalone_rtio_analyzer_fifo_readable = 1'd0;
wire main_genericstandalone_rtio_analyzer_fifo_syncfifo_we;
wire main_genericstandalone_rtio_analyzer_fifo_syncfifo_writable;
wire main_genericstandalone_rtio_analyzer_fifo_syncfifo_re;
wire main_genericstandalone_rtio_analyzer_fifo_syncfifo_readable;
wire [256:0] main_genericstandalone_rtio_analyzer_fifo_syncfifo_din;
wire [256:0] main_genericstandalone_rtio_analyzer_fifo_syncfifo_dout;
reg [7:0] main_genericstandalone_rtio_analyzer_fifo_level0 = 8'd0;
reg main_genericstandalone_rtio_analyzer_fifo_replace = 1'd0;
reg [6:0] main_genericstandalone_rtio_analyzer_fifo_produce = 7'd0;
reg [6:0] main_genericstandalone_rtio_analyzer_fifo_consume = 7'd0;
reg [6:0] main_genericstandalone_rtio_analyzer_fifo_wrport_adr;
wire [256:0] main_genericstandalone_rtio_analyzer_fifo_wrport_dat_r;
wire main_genericstandalone_rtio_analyzer_fifo_wrport_we;
wire [256:0] main_genericstandalone_rtio_analyzer_fifo_wrport_dat_w;
wire main_genericstandalone_rtio_analyzer_fifo_do_read0;
wire [6:0] main_genericstandalone_rtio_analyzer_fifo_rdport_adr;
wire [256:0] main_genericstandalone_rtio_analyzer_fifo_rdport_dat_r;
wire main_genericstandalone_rtio_analyzer_fifo_rdport_re;
wire [7:0] main_genericstandalone_rtio_analyzer_fifo_level1;
wire main_genericstandalone_rtio_analyzer_fifo_almost_full;
wire [255:0] main_genericstandalone_rtio_analyzer_fifo_fifo_in_payload_data;
wire main_genericstandalone_rtio_analyzer_fifo_fifo_in_eop;
wire [255:0] main_genericstandalone_rtio_analyzer_fifo_fifo_out_payload_data;
wire main_genericstandalone_rtio_analyzer_fifo_fifo_out_eop;
reg [5:0] main_genericstandalone_rtio_analyzer_fifo_transfer_count = 6'd63;
wire main_genericstandalone_rtio_analyzer_fifo_transfer_count_ce;
wire main_genericstandalone_rtio_analyzer_fifo_transfer_count_rst;
reg main_genericstandalone_rtio_analyzer_fifo_activated = 1'd0;
reg [7:0] main_genericstandalone_rtio_analyzer_fifo_eop_count = 8'd0;
reg [7:0] main_genericstandalone_rtio_analyzer_fifo_eop_count_next;
wire main_genericstandalone_rtio_analyzer_fifo_has_pending_eop;
wire main_genericstandalone_rtio_analyzer_fifo_do_write;
wire main_genericstandalone_rtio_analyzer_fifo_do_read1;
wire main_genericstandalone_rtio_analyzer_converter_sink_stb;
wire main_genericstandalone_rtio_analyzer_converter_sink_ack;
wire main_genericstandalone_rtio_analyzer_converter_sink_last;
wire main_genericstandalone_rtio_analyzer_converter_sink_eop;
wire [255:0] main_genericstandalone_rtio_analyzer_converter_sink_payload_data;
wire main_genericstandalone_rtio_analyzer_converter_source_stb;
wire main_genericstandalone_rtio_analyzer_converter_source_ack;
wire main_genericstandalone_rtio_analyzer_converter_source_last;
wire main_genericstandalone_rtio_analyzer_converter_source_eop;
reg [127:0] main_genericstandalone_rtio_analyzer_converter_source_payload_data;
wire main_genericstandalone_rtio_analyzer_converter_source_payload_valid_token_count;
reg main_genericstandalone_rtio_analyzer_converter_mux = 1'd0;
wire main_genericstandalone_rtio_analyzer_converter_last;
wire main_genericstandalone_rtio_analyzer_dma_reset_re;
wire main_genericstandalone_rtio_analyzer_dma_reset_r;
reg main_genericstandalone_rtio_analyzer_dma_reset_w = 1'd0;
reg [32:0] main_genericstandalone_rtio_analyzer_dma_base_address_storage_full = 33'd0;
wire [28:0] main_genericstandalone_rtio_analyzer_dma_base_address_storage;
reg main_genericstandalone_rtio_analyzer_dma_base_address_re = 1'd0;
reg [32:0] main_genericstandalone_rtio_analyzer_dma_last_address_storage_full = 33'd0;
wire [28:0] main_genericstandalone_rtio_analyzer_dma_last_address_storage;
reg main_genericstandalone_rtio_analyzer_dma_last_address_re = 1'd0;
wire [63:0] main_genericstandalone_rtio_analyzer_dma_status;
wire main_genericstandalone_rtio_analyzer_dma_sink_stb;
wire main_genericstandalone_rtio_analyzer_dma_sink_ack;
wire main_genericstandalone_rtio_analyzer_dma_sink_last;
wire main_genericstandalone_rtio_analyzer_dma_sink_eop;
wire [127:0] main_genericstandalone_rtio_analyzer_dma_sink_payload_data;
wire main_genericstandalone_rtio_analyzer_dma_sink_payload_valid_token_count;
reg [58:0] main_genericstandalone_rtio_analyzer_dma_message_count = 59'd0;
reg main_genericstandalone_rtio_analyzer_enable_r = 1'd0;
reg [1:0] builder_rtiosyscrg_state = 2'd0;
reg [1:0] builder_rtiosyscrg_next_state;
reg [15:0] main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value0;
reg main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value_ce0;
reg main_genericstandalone_genericstandalone_crg_o_switch_rtiosyscrg_next_value1;
reg main_genericstandalone_genericstandalone_crg_o_switch_rtiosyscrg_next_value_ce1;
reg [5:0] builder_minicon_state = 6'd0;
reg [5:0] builder_minicon_next_state;
reg [2:0] builder_cache_state = 3'd0;
reg [2:0] builder_cache_next_state;
reg builder_icap_state = 1'd0;
reg builder_icap_next_state;
reg [3:0] main_genericstandalone_genericstandalone_icap_counter1_icap_next_value;
reg main_genericstandalone_genericstandalone_icap_counter1_icap_next_value_ce;
reg [2:0] builder_a7_1000basex_transmitpath_state = 3'd0;
reg [2:0] builder_a7_1000basex_transmitpath_next_state;
reg main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value;
reg main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value_ce;
reg [2:0] builder_a7_1000basex_receivepath_state = 3'd0;
reg [2:0] builder_a7_1000basex_receivepath_next_state;
reg [2:0] builder_a7_1000basex_fsm_state = 3'd0;
reg [2:0] builder_a7_1000basex_fsm_next_state;
reg [1:0] builder_a7_1000basex_gtptxinit_state = 2'd0;
reg [1:0] builder_a7_1000basex_gtptxinit_next_state;
reg [3:0] builder_a7_1000basex_gtprxinit_state = 4'd0;
reg [3:0] builder_a7_1000basex_gtprxinit_next_state;
reg [15:0] main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value;
reg main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value_ce;
reg builder_liteethmacgap_state = 1'd0;
reg builder_liteethmacgap_next_state;
reg [1:0] builder_liteethmacpreambleinserter_state = 2'd0;
reg [1:0] builder_liteethmacpreambleinserter_next_state;
reg builder_liteethmacpreamblechecker_state = 1'd0;
reg builder_liteethmacpreamblechecker_next_state;
reg [1:0] builder_liteethmaccrc32inserter_state = 2'd0;
reg [1:0] builder_liteethmaccrc32inserter_next_state;
reg [1:0] builder_liteethmaccrc32checker_state = 2'd0;
reg [1:0] builder_liteethmaccrc32checker_next_state;
reg builder_liteethmacpaddinginserter_state = 1'd0;
reg builder_liteethmacpaddinginserter_next_state;
reg [1:0] builder_liteethmacsramwriter_state = 2'd0;
reg [1:0] builder_liteethmacsramwriter_next_state;
reg [31:0] main_genericstandalone_sram17_status_liteethmac_next_value;
reg main_genericstandalone_sram17_status_liteethmac_next_value_ce;
reg [1:0] builder_liteethmacsramreader_state = 2'd0;
reg [1:0] builder_liteethmacsramreader_next_state;
wire [28:0] builder_shared_adr;
wire [63:0] builder_shared_dat_w;
wire [63:0] builder_shared_dat_r;
wire [7:0] builder_shared_sel;
wire builder_shared_cyc;
wire builder_shared_stb;
wire builder_shared_ack;
wire builder_shared_we;
wire [2:0] builder_shared_cti;
wire [1:0] builder_shared_bte;
wire builder_shared_err;
wire [1:0] builder_request;
reg builder_grant = 1'd0;
reg [4:0] builder_slave_sel;
reg [4:0] builder_slave_sel_r = 5'd0;
reg [2:0] builder_spimaster0_state = 3'd0;
reg [2:0] builder_spimaster0_next_state;
reg builder_ad9910monitor0_state = 1'd0;
reg builder_ad9910monitor0_next_state;
reg [15:0] builder_ad9910monitor0_next_value;
reg builder_ad9910monitor0_next_value_ce;
reg [31:0] main_urukulmonitor0_ftw0_ad9910monitor0_next_value;
reg main_urukulmonitor0_ftw0_ad9910monitor0_next_value_ce;
reg builder_ad9910monitor1_state = 1'd0;
reg builder_ad9910monitor1_next_state;
reg [15:0] builder_ad9910monitor1_next_value;
reg builder_ad9910monitor1_next_value_ce;
reg [31:0] main_urukulmonitor0_ftw1_ad9910monitor1_next_value;
reg main_urukulmonitor0_ftw1_ad9910monitor1_next_value_ce;
reg builder_ad9910monitor2_state = 1'd0;
reg builder_ad9910monitor2_next_state;
reg [15:0] builder_ad9910monitor2_next_value;
reg builder_ad9910monitor2_next_value_ce;
reg [31:0] main_urukulmonitor0_ftw2_ad9910monitor2_next_value;
reg main_urukulmonitor0_ftw2_ad9910monitor2_next_value_ce;
reg builder_ad9910monitor3_state = 1'd0;
reg builder_ad9910monitor3_next_state;
reg [15:0] builder_ad9910monitor3_next_value;
reg builder_ad9910monitor3_next_value_ce;
reg [31:0] main_urukulmonitor0_ftw3_ad9910monitor3_next_value;
reg main_urukulmonitor0_ftw3_ad9910monitor3_next_value_ce;
reg [2:0] builder_spimaster1_state = 3'd0;
reg [2:0] builder_spimaster1_next_state;
reg builder_ad9912monitor0_state = 1'd0;
reg builder_ad9912monitor0_next_state;
reg [15:0] builder_ad9912monitor0_t_next_value;
reg builder_ad9912monitor0_t_next_value_ce;
reg [15:0] builder_ad9912monitor0_f_next_value;
reg builder_ad9912monitor0_f_next_value_ce;
reg builder_ad9912monitor1_state = 1'd0;
reg builder_ad9912monitor1_next_state;
reg [15:0] builder_ad9912monitor1_t_next_value;
reg builder_ad9912monitor1_t_next_value_ce;
reg [15:0] builder_ad9912monitor1_f_next_value;
reg builder_ad9912monitor1_f_next_value_ce;
reg builder_ad9912monitor2_state = 1'd0;
reg builder_ad9912monitor2_next_state;
reg [15:0] builder_ad9912monitor2_t_next_value;
reg builder_ad9912monitor2_t_next_value_ce;
reg [15:0] builder_ad9912monitor2_f_next_value;
reg builder_ad9912monitor2_f_next_value_ce;
reg builder_ad9912monitor3_state = 1'd0;
reg builder_ad9912monitor3_next_state;
reg [15:0] builder_ad9912monitor3_t_next_value;
reg builder_ad9912monitor3_t_next_value_ce;
reg [15:0] builder_ad9912monitor3_f_next_value;
reg builder_ad9912monitor3_f_next_value_ce;
reg [2:0] builder_spimaster2_state = 3'd0;
reg [2:0] builder_spimaster2_next_state;
reg [2:0] builder_spimaster3_state = 3'd0;
reg [2:0] builder_spimaster3_next_state;
reg [2:0] builder_spimaster4_state = 3'd0;
reg [2:0] builder_spimaster4_next_state;
reg [1:0] builder_clockdomainsrenamer_resetinserter_state = 2'd0;
reg [1:0] builder_clockdomainsrenamer_resetinserter_next_state;
reg [1:0] builder_clockdomainsrenamer_recordconverter_state = 2'd0;
reg [1:0] builder_clockdomainsrenamer_recordconverter_next_state;
reg [2:0] builder_clockdomainsrenamer_crimaster_state = 3'd0;
reg [2:0] builder_clockdomainsrenamer_crimaster_next_state;
reg [2:0] builder_clockdomainsrenamer_fsm_state = 3'd0;
reg [2:0] builder_clockdomainsrenamer_fsm_next_state;
wire [1:0] builder_sdram_cpulevel_arbiter_request;
reg builder_sdram_cpulevel_arbiter_grant = 1'd0;
wire [2:0] builder_sdram_native_arbiter_request;
reg [1:0] builder_sdram_native_arbiter_grant = 2'd0;
wire [28:0] builder_genericstandalone_shared_adr;
wire [63:0] builder_genericstandalone_shared_dat_w;
wire [63:0] builder_genericstandalone_shared_dat_r;
wire [7:0] builder_genericstandalone_shared_sel;
wire builder_genericstandalone_shared_cyc;
wire builder_genericstandalone_shared_stb;
wire builder_genericstandalone_shared_ack;
wire builder_genericstandalone_shared_we;
wire [2:0] builder_genericstandalone_shared_cti;
wire [1:0] builder_genericstandalone_shared_bte;
wire builder_genericstandalone_shared_err;
wire [1:0] builder_genericstandalone_request;
reg builder_genericstandalone_grant = 1'd0;
reg [5:0] builder_genericstandalone_slave_sel;
reg [5:0] builder_genericstandalone_slave_sel_r = 6'd0;
wire [13:0] builder_genericstandalone_interface0_bank_bus_adr;
wire builder_genericstandalone_interface0_bank_bus_we;
wire [7:0] builder_genericstandalone_interface0_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface0_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank0_switch_done_re;
wire builder_genericstandalone_csrbank0_switch_done_r;
wire builder_genericstandalone_csrbank0_switch_done_w;
wire builder_genericstandalone_csrbank0_clock_sel0_re;
wire builder_genericstandalone_csrbank0_clock_sel0_r;
wire builder_genericstandalone_csrbank0_clock_sel0_w;
wire builder_genericstandalone_csrbank0_sel;
wire [13:0] builder_genericstandalone_interface1_bank_bus_adr;
wire builder_genericstandalone_interface1_bank_bus_we;
wire [7:0] builder_genericstandalone_interface1_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface1_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank1_dly_sel0_re;
wire [1:0] builder_genericstandalone_csrbank1_dly_sel0_r;
wire [1:0] builder_genericstandalone_csrbank1_dly_sel0_w;
wire builder_genericstandalone_csrbank1_sel;
wire [13:0] builder_genericstandalone_interface2_bank_bus_adr;
wire builder_genericstandalone_interface2_bank_bus_we;
wire [7:0] builder_genericstandalone_interface2_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface2_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank2_control0_re;
wire [3:0] builder_genericstandalone_csrbank2_control0_r;
wire [3:0] builder_genericstandalone_csrbank2_control0_w;
wire builder_genericstandalone_csrbank2_pi0_command0_re;
wire [5:0] builder_genericstandalone_csrbank2_pi0_command0_r;
wire [5:0] builder_genericstandalone_csrbank2_pi0_command0_w;
wire builder_genericstandalone_csrbank2_pi0_address1_re;
wire [6:0] builder_genericstandalone_csrbank2_pi0_address1_r;
wire [6:0] builder_genericstandalone_csrbank2_pi0_address1_w;
wire builder_genericstandalone_csrbank2_pi0_address0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_address0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_address0_w;
wire builder_genericstandalone_csrbank2_pi0_baddress0_re;
wire [2:0] builder_genericstandalone_csrbank2_pi0_baddress0_r;
wire [2:0] builder_genericstandalone_csrbank2_pi0_baddress0_w;
wire builder_genericstandalone_csrbank2_pi0_wrdata3_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_wrdata3_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_wrdata3_w;
wire builder_genericstandalone_csrbank2_pi0_wrdata2_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_wrdata2_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_wrdata2_w;
wire builder_genericstandalone_csrbank2_pi0_wrdata1_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_wrdata1_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_wrdata1_w;
wire builder_genericstandalone_csrbank2_pi0_wrdata0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_wrdata0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_wrdata0_w;
wire builder_genericstandalone_csrbank2_pi0_rddata3_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_rddata3_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_rddata3_w;
wire builder_genericstandalone_csrbank2_pi0_rddata2_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_rddata2_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_rddata2_w;
wire builder_genericstandalone_csrbank2_pi0_rddata1_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_rddata1_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_rddata1_w;
wire builder_genericstandalone_csrbank2_pi0_rddata0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi0_rddata0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi0_rddata0_w;
wire builder_genericstandalone_csrbank2_pi1_command0_re;
wire [5:0] builder_genericstandalone_csrbank2_pi1_command0_r;
wire [5:0] builder_genericstandalone_csrbank2_pi1_command0_w;
wire builder_genericstandalone_csrbank2_pi1_address1_re;
wire [6:0] builder_genericstandalone_csrbank2_pi1_address1_r;
wire [6:0] builder_genericstandalone_csrbank2_pi1_address1_w;
wire builder_genericstandalone_csrbank2_pi1_address0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_address0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_address0_w;
wire builder_genericstandalone_csrbank2_pi1_baddress0_re;
wire [2:0] builder_genericstandalone_csrbank2_pi1_baddress0_r;
wire [2:0] builder_genericstandalone_csrbank2_pi1_baddress0_w;
wire builder_genericstandalone_csrbank2_pi1_wrdata3_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_wrdata3_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_wrdata3_w;
wire builder_genericstandalone_csrbank2_pi1_wrdata2_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_wrdata2_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_wrdata2_w;
wire builder_genericstandalone_csrbank2_pi1_wrdata1_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_wrdata1_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_wrdata1_w;
wire builder_genericstandalone_csrbank2_pi1_wrdata0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_wrdata0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_wrdata0_w;
wire builder_genericstandalone_csrbank2_pi1_rddata3_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_rddata3_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_rddata3_w;
wire builder_genericstandalone_csrbank2_pi1_rddata2_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_rddata2_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_rddata2_w;
wire builder_genericstandalone_csrbank2_pi1_rddata1_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_rddata1_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_rddata1_w;
wire builder_genericstandalone_csrbank2_pi1_rddata0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi1_rddata0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi1_rddata0_w;
wire builder_genericstandalone_csrbank2_pi2_command0_re;
wire [5:0] builder_genericstandalone_csrbank2_pi2_command0_r;
wire [5:0] builder_genericstandalone_csrbank2_pi2_command0_w;
wire builder_genericstandalone_csrbank2_pi2_address1_re;
wire [6:0] builder_genericstandalone_csrbank2_pi2_address1_r;
wire [6:0] builder_genericstandalone_csrbank2_pi2_address1_w;
wire builder_genericstandalone_csrbank2_pi2_address0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_address0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_address0_w;
wire builder_genericstandalone_csrbank2_pi2_baddress0_re;
wire [2:0] builder_genericstandalone_csrbank2_pi2_baddress0_r;
wire [2:0] builder_genericstandalone_csrbank2_pi2_baddress0_w;
wire builder_genericstandalone_csrbank2_pi2_wrdata3_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_wrdata3_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_wrdata3_w;
wire builder_genericstandalone_csrbank2_pi2_wrdata2_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_wrdata2_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_wrdata2_w;
wire builder_genericstandalone_csrbank2_pi2_wrdata1_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_wrdata1_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_wrdata1_w;
wire builder_genericstandalone_csrbank2_pi2_wrdata0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_wrdata0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_wrdata0_w;
wire builder_genericstandalone_csrbank2_pi2_rddata3_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_rddata3_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_rddata3_w;
wire builder_genericstandalone_csrbank2_pi2_rddata2_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_rddata2_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_rddata2_w;
wire builder_genericstandalone_csrbank2_pi2_rddata1_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_rddata1_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_rddata1_w;
wire builder_genericstandalone_csrbank2_pi2_rddata0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi2_rddata0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi2_rddata0_w;
wire builder_genericstandalone_csrbank2_pi3_command0_re;
wire [5:0] builder_genericstandalone_csrbank2_pi3_command0_r;
wire [5:0] builder_genericstandalone_csrbank2_pi3_command0_w;
wire builder_genericstandalone_csrbank2_pi3_address1_re;
wire [6:0] builder_genericstandalone_csrbank2_pi3_address1_r;
wire [6:0] builder_genericstandalone_csrbank2_pi3_address1_w;
wire builder_genericstandalone_csrbank2_pi3_address0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_address0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_address0_w;
wire builder_genericstandalone_csrbank2_pi3_baddress0_re;
wire [2:0] builder_genericstandalone_csrbank2_pi3_baddress0_r;
wire [2:0] builder_genericstandalone_csrbank2_pi3_baddress0_w;
wire builder_genericstandalone_csrbank2_pi3_wrdata3_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_wrdata3_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_wrdata3_w;
wire builder_genericstandalone_csrbank2_pi3_wrdata2_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_wrdata2_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_wrdata2_w;
wire builder_genericstandalone_csrbank2_pi3_wrdata1_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_wrdata1_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_wrdata1_w;
wire builder_genericstandalone_csrbank2_pi3_wrdata0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_wrdata0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_wrdata0_w;
wire builder_genericstandalone_csrbank2_pi3_rddata3_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_rddata3_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_rddata3_w;
wire builder_genericstandalone_csrbank2_pi3_rddata2_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_rddata2_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_rddata2_w;
wire builder_genericstandalone_csrbank2_pi3_rddata1_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_rddata1_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_rddata1_w;
wire builder_genericstandalone_csrbank2_pi3_rddata0_re;
wire [7:0] builder_genericstandalone_csrbank2_pi3_rddata0_r;
wire [7:0] builder_genericstandalone_csrbank2_pi3_rddata0_w;
wire builder_genericstandalone_csrbank2_sel;
wire [13:0] builder_genericstandalone_interface3_bank_bus_adr;
wire builder_genericstandalone_interface3_bank_bus_we;
wire [7:0] builder_genericstandalone_interface3_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface3_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank3_out0_re;
wire builder_genericstandalone_csrbank3_out0_r;
wire builder_genericstandalone_csrbank3_out0_w;
wire builder_genericstandalone_csrbank3_sel;
wire [13:0] builder_genericstandalone_interface4_bank_bus_adr;
wire builder_genericstandalone_interface4_bank_bus_we;
wire [7:0] builder_genericstandalone_interface4_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface4_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank4_sram_writer_slot_re;
wire [1:0] builder_genericstandalone_csrbank4_sram_writer_slot_r;
wire [1:0] builder_genericstandalone_csrbank4_sram_writer_slot_w;
wire builder_genericstandalone_csrbank4_sram_writer_length1_re;
wire [2:0] builder_genericstandalone_csrbank4_sram_writer_length1_r;
wire [2:0] builder_genericstandalone_csrbank4_sram_writer_length1_w;
wire builder_genericstandalone_csrbank4_sram_writer_length0_re;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_length0_r;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_length0_w;
wire builder_genericstandalone_csrbank4_sram_writer_errors3_re;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_errors3_r;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_errors3_w;
wire builder_genericstandalone_csrbank4_sram_writer_errors2_re;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_errors2_r;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_errors2_w;
wire builder_genericstandalone_csrbank4_sram_writer_errors1_re;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_errors1_r;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_errors1_w;
wire builder_genericstandalone_csrbank4_sram_writer_errors0_re;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_errors0_r;
wire [7:0] builder_genericstandalone_csrbank4_sram_writer_errors0_w;
wire builder_genericstandalone_csrbank4_sram_writer_ev_enable0_re;
wire builder_genericstandalone_csrbank4_sram_writer_ev_enable0_r;
wire builder_genericstandalone_csrbank4_sram_writer_ev_enable0_w;
wire builder_genericstandalone_csrbank4_sram_reader_ready_re;
wire builder_genericstandalone_csrbank4_sram_reader_ready_r;
wire builder_genericstandalone_csrbank4_sram_reader_ready_w;
wire builder_genericstandalone_csrbank4_sram_reader_slot0_re;
wire [1:0] builder_genericstandalone_csrbank4_sram_reader_slot0_r;
wire [1:0] builder_genericstandalone_csrbank4_sram_reader_slot0_w;
wire builder_genericstandalone_csrbank4_sram_reader_length1_re;
wire [2:0] builder_genericstandalone_csrbank4_sram_reader_length1_r;
wire [2:0] builder_genericstandalone_csrbank4_sram_reader_length1_w;
wire builder_genericstandalone_csrbank4_sram_reader_length0_re;
wire [7:0] builder_genericstandalone_csrbank4_sram_reader_length0_r;
wire [7:0] builder_genericstandalone_csrbank4_sram_reader_length0_w;
wire builder_genericstandalone_csrbank4_sram_reader_ev_enable0_re;
wire builder_genericstandalone_csrbank4_sram_reader_ev_enable0_r;
wire builder_genericstandalone_csrbank4_sram_reader_ev_enable0_w;
wire builder_genericstandalone_csrbank4_preamble_errors3_re;
wire [7:0] builder_genericstandalone_csrbank4_preamble_errors3_r;
wire [7:0] builder_genericstandalone_csrbank4_preamble_errors3_w;
wire builder_genericstandalone_csrbank4_preamble_errors2_re;
wire [7:0] builder_genericstandalone_csrbank4_preamble_errors2_r;
wire [7:0] builder_genericstandalone_csrbank4_preamble_errors2_w;
wire builder_genericstandalone_csrbank4_preamble_errors1_re;
wire [7:0] builder_genericstandalone_csrbank4_preamble_errors1_r;
wire [7:0] builder_genericstandalone_csrbank4_preamble_errors1_w;
wire builder_genericstandalone_csrbank4_preamble_errors0_re;
wire [7:0] builder_genericstandalone_csrbank4_preamble_errors0_r;
wire [7:0] builder_genericstandalone_csrbank4_preamble_errors0_w;
wire builder_genericstandalone_csrbank4_crc_errors3_re;
wire [7:0] builder_genericstandalone_csrbank4_crc_errors3_r;
wire [7:0] builder_genericstandalone_csrbank4_crc_errors3_w;
wire builder_genericstandalone_csrbank4_crc_errors2_re;
wire [7:0] builder_genericstandalone_csrbank4_crc_errors2_r;
wire [7:0] builder_genericstandalone_csrbank4_crc_errors2_w;
wire builder_genericstandalone_csrbank4_crc_errors1_re;
wire [7:0] builder_genericstandalone_csrbank4_crc_errors1_r;
wire [7:0] builder_genericstandalone_csrbank4_crc_errors1_w;
wire builder_genericstandalone_csrbank4_crc_errors0_re;
wire [7:0] builder_genericstandalone_csrbank4_crc_errors0_r;
wire [7:0] builder_genericstandalone_csrbank4_crc_errors0_w;
wire builder_genericstandalone_csrbank4_sel;
wire [13:0] builder_genericstandalone_interface5_bank_bus_adr;
wire builder_genericstandalone_interface5_bank_bus_we;
wire [7:0] builder_genericstandalone_interface5_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface5_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank5_in_re;
wire [1:0] builder_genericstandalone_csrbank5_in_r;
wire [1:0] builder_genericstandalone_csrbank5_in_w;
wire builder_genericstandalone_csrbank5_out0_re;
wire [1:0] builder_genericstandalone_csrbank5_out0_r;
wire [1:0] builder_genericstandalone_csrbank5_out0_w;
wire builder_genericstandalone_csrbank5_oe0_re;
wire [1:0] builder_genericstandalone_csrbank5_oe0_r;
wire [1:0] builder_genericstandalone_csrbank5_oe0_w;
wire builder_genericstandalone_csrbank5_sel;
wire [13:0] builder_genericstandalone_interface6_bank_bus_adr;
wire builder_genericstandalone_interface6_bank_bus_we;
wire [7:0] builder_genericstandalone_interface6_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface6_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank6_sel;
wire [13:0] builder_genericstandalone_interface7_bank_bus_adr;
wire builder_genericstandalone_interface7_bank_bus_we;
wire [7:0] builder_genericstandalone_interface7_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface7_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank7_address0_re;
wire [7:0] builder_genericstandalone_csrbank7_address0_r;
wire [7:0] builder_genericstandalone_csrbank7_address0_w;
wire builder_genericstandalone_csrbank7_data_re;
wire [7:0] builder_genericstandalone_csrbank7_data_r;
wire [7:0] builder_genericstandalone_csrbank7_data_w;
wire builder_genericstandalone_csrbank7_sel;
wire [13:0] builder_genericstandalone_interface8_bank_bus_adr;
wire builder_genericstandalone_interface8_bank_bus_we;
wire [7:0] builder_genericstandalone_interface8_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface8_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank8_reset0_re;
wire builder_genericstandalone_csrbank8_reset0_r;
wire builder_genericstandalone_csrbank8_reset0_w;
wire builder_genericstandalone_csrbank8_sel;
wire [13:0] builder_genericstandalone_interface9_bank_bus_adr;
wire builder_genericstandalone_interface9_bank_bus_we;
wire [7:0] builder_genericstandalone_interface9_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface9_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank9_enable0_re;
wire builder_genericstandalone_csrbank9_enable0_r;
wire builder_genericstandalone_csrbank9_enable0_w;
wire builder_genericstandalone_csrbank9_busy_re;
wire builder_genericstandalone_csrbank9_busy_r;
wire builder_genericstandalone_csrbank9_busy_w;
wire builder_genericstandalone_csrbank9_message_encoder_overflow_re;
wire builder_genericstandalone_csrbank9_message_encoder_overflow_r;
wire builder_genericstandalone_csrbank9_message_encoder_overflow_w;
wire builder_genericstandalone_csrbank9_dma_base_address4_re;
wire builder_genericstandalone_csrbank9_dma_base_address4_r;
wire builder_genericstandalone_csrbank9_dma_base_address4_w;
wire builder_genericstandalone_csrbank9_dma_base_address3_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_base_address3_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_base_address3_w;
wire builder_genericstandalone_csrbank9_dma_base_address2_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_base_address2_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_base_address2_w;
wire builder_genericstandalone_csrbank9_dma_base_address1_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_base_address1_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_base_address1_w;
wire builder_genericstandalone_csrbank9_dma_base_address0_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_base_address0_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_base_address0_w;
wire builder_genericstandalone_csrbank9_dma_last_address4_re;
wire builder_genericstandalone_csrbank9_dma_last_address4_r;
wire builder_genericstandalone_csrbank9_dma_last_address4_w;
wire builder_genericstandalone_csrbank9_dma_last_address3_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_last_address3_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_last_address3_w;
wire builder_genericstandalone_csrbank9_dma_last_address2_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_last_address2_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_last_address2_w;
wire builder_genericstandalone_csrbank9_dma_last_address1_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_last_address1_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_last_address1_w;
wire builder_genericstandalone_csrbank9_dma_last_address0_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_last_address0_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_last_address0_w;
wire builder_genericstandalone_csrbank9_dma_byte_count7_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count7_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count7_w;
wire builder_genericstandalone_csrbank9_dma_byte_count6_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count6_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count6_w;
wire builder_genericstandalone_csrbank9_dma_byte_count5_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count5_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count5_w;
wire builder_genericstandalone_csrbank9_dma_byte_count4_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count4_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count4_w;
wire builder_genericstandalone_csrbank9_dma_byte_count3_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count3_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count3_w;
wire builder_genericstandalone_csrbank9_dma_byte_count2_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count2_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count2_w;
wire builder_genericstandalone_csrbank9_dma_byte_count1_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count1_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count1_w;
wire builder_genericstandalone_csrbank9_dma_byte_count0_re;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count0_r;
wire [7:0] builder_genericstandalone_csrbank9_dma_byte_count0_w;
wire builder_genericstandalone_csrbank9_sel;
wire [13:0] builder_genericstandalone_interface10_bank_bus_adr;
wire builder_genericstandalone_interface10_bank_bus_we;
wire [7:0] builder_genericstandalone_interface10_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface10_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank10_sed_spread_enable0_re;
wire builder_genericstandalone_csrbank10_sed_spread_enable0_r;
wire builder_genericstandalone_csrbank10_sed_spread_enable0_w;
wire builder_genericstandalone_csrbank10_collision_channel1_re;
wire [7:0] builder_genericstandalone_csrbank10_collision_channel1_r;
wire [7:0] builder_genericstandalone_csrbank10_collision_channel1_w;
wire builder_genericstandalone_csrbank10_collision_channel0_re;
wire [7:0] builder_genericstandalone_csrbank10_collision_channel0_r;
wire [7:0] builder_genericstandalone_csrbank10_collision_channel0_w;
wire builder_genericstandalone_csrbank10_busy_channel1_re;
wire [7:0] builder_genericstandalone_csrbank10_busy_channel1_r;
wire [7:0] builder_genericstandalone_csrbank10_busy_channel1_w;
wire builder_genericstandalone_csrbank10_busy_channel0_re;
wire [7:0] builder_genericstandalone_csrbank10_busy_channel0_r;
wire [7:0] builder_genericstandalone_csrbank10_busy_channel0_w;
wire builder_genericstandalone_csrbank10_sequence_error_channel1_re;
wire [7:0] builder_genericstandalone_csrbank10_sequence_error_channel1_r;
wire [7:0] builder_genericstandalone_csrbank10_sequence_error_channel1_w;
wire builder_genericstandalone_csrbank10_sequence_error_channel0_re;
wire [7:0] builder_genericstandalone_csrbank10_sequence_error_channel0_r;
wire [7:0] builder_genericstandalone_csrbank10_sequence_error_channel0_w;
wire builder_genericstandalone_csrbank10_sel;
wire [13:0] builder_genericstandalone_interface11_bank_bus_adr;
wire builder_genericstandalone_interface11_bank_bus_we;
wire [7:0] builder_genericstandalone_interface11_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface11_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank11_mon_chan_sel0_re;
wire [5:0] builder_genericstandalone_csrbank11_mon_chan_sel0_r;
wire [5:0] builder_genericstandalone_csrbank11_mon_chan_sel0_w;
wire builder_genericstandalone_csrbank11_mon_probe_sel0_re;
wire [4:0] builder_genericstandalone_csrbank11_mon_probe_sel0_r;
wire [4:0] builder_genericstandalone_csrbank11_mon_probe_sel0_w;
wire builder_genericstandalone_csrbank11_mon_value3_re;
wire [7:0] builder_genericstandalone_csrbank11_mon_value3_r;
wire [7:0] builder_genericstandalone_csrbank11_mon_value3_w;
wire builder_genericstandalone_csrbank11_mon_value2_re;
wire [7:0] builder_genericstandalone_csrbank11_mon_value2_r;
wire [7:0] builder_genericstandalone_csrbank11_mon_value2_w;
wire builder_genericstandalone_csrbank11_mon_value1_re;
wire [7:0] builder_genericstandalone_csrbank11_mon_value1_r;
wire [7:0] builder_genericstandalone_csrbank11_mon_value1_w;
wire builder_genericstandalone_csrbank11_mon_value0_re;
wire [7:0] builder_genericstandalone_csrbank11_mon_value0_r;
wire [7:0] builder_genericstandalone_csrbank11_mon_value0_w;
wire builder_genericstandalone_csrbank11_inj_chan_sel0_re;
wire [5:0] builder_genericstandalone_csrbank11_inj_chan_sel0_r;
wire [5:0] builder_genericstandalone_csrbank11_inj_chan_sel0_w;
wire builder_genericstandalone_csrbank11_inj_override_sel0_re;
wire [1:0] builder_genericstandalone_csrbank11_inj_override_sel0_r;
wire [1:0] builder_genericstandalone_csrbank11_inj_override_sel0_w;
wire builder_genericstandalone_csrbank11_sel;
wire [13:0] builder_genericstandalone_interface12_bank_bus_adr;
wire builder_genericstandalone_interface12_bank_bus_we;
wire [7:0] builder_genericstandalone_interface12_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface12_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank12_bitbang0_re;
wire [3:0] builder_genericstandalone_csrbank12_bitbang0_r;
wire [3:0] builder_genericstandalone_csrbank12_bitbang0_w;
wire builder_genericstandalone_csrbank12_miso_re;
wire builder_genericstandalone_csrbank12_miso_r;
wire builder_genericstandalone_csrbank12_miso_w;
wire builder_genericstandalone_csrbank12_bitbang_en0_re;
wire builder_genericstandalone_csrbank12_bitbang_en0_r;
wire builder_genericstandalone_csrbank12_bitbang_en0_w;
wire builder_genericstandalone_csrbank12_sel;
wire [13:0] builder_genericstandalone_interface13_bank_bus_adr;
wire builder_genericstandalone_interface13_bank_bus_we;
wire [7:0] builder_genericstandalone_interface13_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface13_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank13_load7_re;
wire [7:0] builder_genericstandalone_csrbank13_load7_r;
wire [7:0] builder_genericstandalone_csrbank13_load7_w;
wire builder_genericstandalone_csrbank13_load6_re;
wire [7:0] builder_genericstandalone_csrbank13_load6_r;
wire [7:0] builder_genericstandalone_csrbank13_load6_w;
wire builder_genericstandalone_csrbank13_load5_re;
wire [7:0] builder_genericstandalone_csrbank13_load5_r;
wire [7:0] builder_genericstandalone_csrbank13_load5_w;
wire builder_genericstandalone_csrbank13_load4_re;
wire [7:0] builder_genericstandalone_csrbank13_load4_r;
wire [7:0] builder_genericstandalone_csrbank13_load4_w;
wire builder_genericstandalone_csrbank13_load3_re;
wire [7:0] builder_genericstandalone_csrbank13_load3_r;
wire [7:0] builder_genericstandalone_csrbank13_load3_w;
wire builder_genericstandalone_csrbank13_load2_re;
wire [7:0] builder_genericstandalone_csrbank13_load2_r;
wire [7:0] builder_genericstandalone_csrbank13_load2_w;
wire builder_genericstandalone_csrbank13_load1_re;
wire [7:0] builder_genericstandalone_csrbank13_load1_r;
wire [7:0] builder_genericstandalone_csrbank13_load1_w;
wire builder_genericstandalone_csrbank13_load0_re;
wire [7:0] builder_genericstandalone_csrbank13_load0_r;
wire [7:0] builder_genericstandalone_csrbank13_load0_w;
wire builder_genericstandalone_csrbank13_reload7_re;
wire [7:0] builder_genericstandalone_csrbank13_reload7_r;
wire [7:0] builder_genericstandalone_csrbank13_reload7_w;
wire builder_genericstandalone_csrbank13_reload6_re;
wire [7:0] builder_genericstandalone_csrbank13_reload6_r;
wire [7:0] builder_genericstandalone_csrbank13_reload6_w;
wire builder_genericstandalone_csrbank13_reload5_re;
wire [7:0] builder_genericstandalone_csrbank13_reload5_r;
wire [7:0] builder_genericstandalone_csrbank13_reload5_w;
wire builder_genericstandalone_csrbank13_reload4_re;
wire [7:0] builder_genericstandalone_csrbank13_reload4_r;
wire [7:0] builder_genericstandalone_csrbank13_reload4_w;
wire builder_genericstandalone_csrbank13_reload3_re;
wire [7:0] builder_genericstandalone_csrbank13_reload3_r;
wire [7:0] builder_genericstandalone_csrbank13_reload3_w;
wire builder_genericstandalone_csrbank13_reload2_re;
wire [7:0] builder_genericstandalone_csrbank13_reload2_r;
wire [7:0] builder_genericstandalone_csrbank13_reload2_w;
wire builder_genericstandalone_csrbank13_reload1_re;
wire [7:0] builder_genericstandalone_csrbank13_reload1_r;
wire [7:0] builder_genericstandalone_csrbank13_reload1_w;
wire builder_genericstandalone_csrbank13_reload0_re;
wire [7:0] builder_genericstandalone_csrbank13_reload0_r;
wire [7:0] builder_genericstandalone_csrbank13_reload0_w;
wire builder_genericstandalone_csrbank13_en0_re;
wire builder_genericstandalone_csrbank13_en0_r;
wire builder_genericstandalone_csrbank13_en0_w;
wire builder_genericstandalone_csrbank13_value7_re;
wire [7:0] builder_genericstandalone_csrbank13_value7_r;
wire [7:0] builder_genericstandalone_csrbank13_value7_w;
wire builder_genericstandalone_csrbank13_value6_re;
wire [7:0] builder_genericstandalone_csrbank13_value6_r;
wire [7:0] builder_genericstandalone_csrbank13_value6_w;
wire builder_genericstandalone_csrbank13_value5_re;
wire [7:0] builder_genericstandalone_csrbank13_value5_r;
wire [7:0] builder_genericstandalone_csrbank13_value5_w;
wire builder_genericstandalone_csrbank13_value4_re;
wire [7:0] builder_genericstandalone_csrbank13_value4_r;
wire [7:0] builder_genericstandalone_csrbank13_value4_w;
wire builder_genericstandalone_csrbank13_value3_re;
wire [7:0] builder_genericstandalone_csrbank13_value3_r;
wire [7:0] builder_genericstandalone_csrbank13_value3_w;
wire builder_genericstandalone_csrbank13_value2_re;
wire [7:0] builder_genericstandalone_csrbank13_value2_r;
wire [7:0] builder_genericstandalone_csrbank13_value2_w;
wire builder_genericstandalone_csrbank13_value1_re;
wire [7:0] builder_genericstandalone_csrbank13_value1_r;
wire [7:0] builder_genericstandalone_csrbank13_value1_w;
wire builder_genericstandalone_csrbank13_value0_re;
wire [7:0] builder_genericstandalone_csrbank13_value0_r;
wire [7:0] builder_genericstandalone_csrbank13_value0_w;
wire builder_genericstandalone_csrbank13_ev_enable0_re;
wire builder_genericstandalone_csrbank13_ev_enable0_r;
wire builder_genericstandalone_csrbank13_ev_enable0_w;
wire builder_genericstandalone_csrbank13_sel;
wire [13:0] builder_genericstandalone_interface14_bank_bus_adr;
wire builder_genericstandalone_interface14_bank_bus_we;
wire [7:0] builder_genericstandalone_interface14_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface14_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank14_txfull_re;
wire builder_genericstandalone_csrbank14_txfull_r;
wire builder_genericstandalone_csrbank14_txfull_w;
wire builder_genericstandalone_csrbank14_rxempty_re;
wire builder_genericstandalone_csrbank14_rxempty_r;
wire builder_genericstandalone_csrbank14_rxempty_w;
wire builder_genericstandalone_csrbank14_ev_enable0_re;
wire [1:0] builder_genericstandalone_csrbank14_ev_enable0_r;
wire [1:0] builder_genericstandalone_csrbank14_ev_enable0_w;
wire builder_genericstandalone_csrbank14_sel;
wire [13:0] builder_genericstandalone_interface15_bank_bus_adr;
wire builder_genericstandalone_interface15_bank_bus_we;
wire [7:0] builder_genericstandalone_interface15_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface15_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank15_tuning_word3_re;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word3_r;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word3_w;
wire builder_genericstandalone_csrbank15_tuning_word2_re;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word2_r;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word2_w;
wire builder_genericstandalone_csrbank15_tuning_word1_re;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word1_r;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word1_w;
wire builder_genericstandalone_csrbank15_tuning_word0_re;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word0_r;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word0_w;
wire builder_genericstandalone_csrbank15_sel;
wire [13:0] builder_genericstandalone_interface16_bank_bus_adr;
wire builder_genericstandalone_interface16_bank_bus_we;
wire [7:0] builder_genericstandalone_interface16_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface16_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank16_status_re;
wire [7:0] builder_genericstandalone_csrbank16_status_r;
wire [7:0] builder_genericstandalone_csrbank16_status_w;
wire builder_genericstandalone_csrbank16_sel;
wire [63:0] builder_slice_proxy0;
wire [63:0] builder_slice_proxy1;
wire [63:0] builder_slice_proxy2;
wire [63:0] builder_slice_proxy3;
wire [63:0] builder_slice_proxy4;
wire [63:0] builder_slice_proxy5;
wire [63:0] builder_slice_proxy6;
wire [63:0] builder_slice_proxy7;
wire [63:0] builder_slice_proxy8;
wire [63:0] builder_slice_proxy9;
wire [63:0] builder_slice_proxy10;
wire [63:0] builder_slice_proxy11;
wire [63:0] builder_slice_proxy12;
wire [63:0] builder_slice_proxy13;
wire [63:0] builder_slice_proxy14;
wire [63:0] builder_slice_proxy15;
wire [63:0] builder_slice_proxy16;
wire [63:0] builder_slice_proxy17;
wire [63:0] builder_slice_proxy18;
wire [63:0] builder_slice_proxy19;
wire [63:0] builder_slice_proxy20;
wire [63:0] builder_slice_proxy21;
wire [63:0] builder_slice_proxy22;
wire [63:0] builder_slice_proxy23;
wire [63:0] builder_slice_proxy24;
wire [63:0] builder_slice_proxy25;
wire [63:0] builder_slice_proxy26;
wire [63:0] builder_slice_proxy27;
wire [63:0] builder_slice_proxy28;
wire [63:0] builder_slice_proxy29;
wire [63:0] builder_slice_proxy30;
wire [63:0] builder_slice_proxy31;
reg [31:0] builder_comb_basiclowerer_self;
reg [28:0] builder_comb_rhs_self0;
reg [63:0] builder_comb_rhs_self1;
reg [7:0] builder_comb_rhs_self2;
reg builder_comb_rhs_self3;
reg builder_comb_rhs_self4;
reg builder_comb_rhs_self5;
reg [2:0] builder_comb_rhs_self6;
reg [1:0] builder_comb_rhs_self7;
wire builder_comb_lhs_self;
reg builder_comb_rhs_self8;
reg builder_comb_rhs_self9;
reg [1:0] builder_comb_rhs_self10;
reg [1:0] builder_comb_rhs_self11;
reg [23:0] builder_comb_rhs_self12;
reg [63:0] builder_comb_rhs_self13;
reg [511:0] builder_comb_rhs_self14;
reg [7:0] builder_comb_rhs_self15;
reg [63:0] builder_comb_rhs_self16;
reg builder_comb_rhs_self17;
reg builder_comb_rhs_self18;
reg builder_comb_rhs_self19;
reg builder_comb_rhs_self20;
reg builder_comb_rhs_self21;
reg builder_comb_rhs_self22;
reg builder_comb_rhs_self23;
reg builder_comb_rhs_self24;
reg builder_comb_rhs_self25;
reg builder_comb_rhs_self26;
reg builder_comb_rhs_self27;
reg builder_comb_rhs_self28;
reg builder_comb_rhs_self29;
reg builder_comb_rhs_self30;
reg builder_comb_rhs_self31;
reg builder_comb_rhs_self32;
reg builder_comb_rhs_self33;
reg builder_comb_rhs_self34;
reg builder_comb_rhs_self35;
reg builder_comb_rhs_self36;
reg builder_comb_rhs_self37;
reg builder_comb_rhs_self38;
reg builder_comb_rhs_self39;
reg builder_comb_rhs_self40;
reg builder_comb_rhs_self41;
reg builder_comb_rhs_self42;
reg builder_comb_rhs_self43;
reg builder_comb_rhs_self44;
reg builder_comb_rhs_self45;
reg builder_comb_rhs_self46;
reg builder_comb_rhs_self47;
reg builder_comb_rhs_self48;
reg builder_comb_rhs_self49;
reg builder_comb_rhs_self50;
reg builder_comb_rhs_self51;
reg builder_comb_rhs_self52;
reg builder_comb_rhs_self53;
reg builder_comb_rhs_self54;
reg builder_comb_rhs_self55;
reg [28:0] builder_comb_rhs_self56;
reg [63:0] builder_comb_rhs_self57;
reg [7:0] builder_comb_rhs_self58;
reg builder_comb_rhs_self59;
reg builder_comb_rhs_self60;
reg builder_comb_rhs_self61;
reg [2:0] builder_comb_rhs_self62;
reg [1:0] builder_comb_rhs_self63;
reg [28:0] builder_comb_rhs_self64;
reg [127:0] builder_comb_rhs_self65;
reg [15:0] builder_comb_rhs_self66;
reg builder_comb_rhs_self67;
reg builder_comb_rhs_self68;
reg builder_comb_rhs_self69;
reg [2:0] builder_comb_rhs_self70;
reg [1:0] builder_comb_rhs_self71;
reg [28:0] builder_comb_rhs_self72;
reg [63:0] builder_comb_rhs_self73;
reg [7:0] builder_comb_rhs_self74;
reg builder_comb_rhs_self75;
reg builder_comb_rhs_self76;
reg builder_comb_rhs_self77;
reg [2:0] builder_comb_rhs_self78;
reg [1:0] builder_comb_rhs_self79;
reg [2:0] builder_sync_t_rhs_self0;
reg [2:0] builder_sync_f_t_self0;
reg [2:0] builder_sync_f_rhs_self0;
reg [4:0] builder_sync_rhs_self0;
reg [5:0] builder_sync_f_rhs_self1;
reg builder_sync_f_rhs_self2;
reg builder_sync_f_rhs_self3;
reg [3:0] builder_sync_rhs_self1;
reg builder_sync_rhs_self2;
reg builder_sync_f_rhs_self4;
reg [60:0] builder_sync_rhs_self3;
reg [60:0] builder_sync_rhs_self4;
reg [60:0] builder_sync_t_lhs_self = 61'd0;
reg builder_sync_basiclowerer_self0;
reg builder_sync_basiclowerer_self1;
reg builder_sync_basiclowerer_self2;
reg builder_sync_basiclowerer_self3;
reg builder_sync_basiclowerer_self4;
reg builder_sync_basiclowerer_self5;
reg builder_sync_basiclowerer_self6;
reg builder_sync_basiclowerer_self7;
reg builder_sync_basiclowerer_self8;
reg builder_sync_basiclowerer_self9;
reg builder_sync_basiclowerer_self10;
reg builder_sync_basiclowerer_self11;
reg builder_sync_basiclowerer_self12;
reg builder_sync_basiclowerer_self13;
reg builder_sync_basiclowerer_self14;
reg builder_sync_basiclowerer_self15;
reg [31:0] builder_sync_t_rhs_self1;
reg [64:0] builder_sync_t_rhs_self2;
reg [7:0] builder_sync_f_t_self1;
reg [6:0] builder_sync_f_t_self2;
reg [7:0] builder_sync_f_t_self3;
reg [6:0] builder_sync_f_t_self4;
reg [7:0] builder_sync_f_t_self5;
reg [6:0] builder_sync_f_t_self6;
reg [7:0] builder_sync_f_t_self7;
reg [6:0] builder_sync_f_t_self8;
reg [7:0] builder_sync_f_t_self9;
reg [6:0] builder_sync_f_t_self10;
reg [7:0] builder_sync_f_t_self11;
reg [6:0] builder_sync_f_t_self12;
reg [7:0] builder_sync_f_t_self13;
reg [6:0] builder_sync_f_t_self14;
reg [7:0] builder_sync_f_t_self15;
reg [6:0] builder_sync_f_t_self16;
reg [7:0] builder_sync_f_t_self17;
reg [6:0] builder_sync_f_t_self18;
reg [7:0] builder_sync_f_t_self19;
reg [6:0] builder_sync_f_t_self20;
reg [7:0] builder_sync_f_t_self21;
reg [6:0] builder_sync_f_t_self22;
reg [7:0] builder_sync_f_t_self23;
reg [6:0] builder_sync_f_t_self24;
reg [7:0] builder_sync_f_t_self25;
reg [6:0] builder_sync_f_t_self26;
reg [7:0] builder_sync_f_t_self27;
reg [6:0] builder_sync_f_t_self28;
reg [7:0] builder_sync_f_t_self29;
reg [6:0] builder_sync_f_t_self30;
reg [7:0] builder_sync_f_t_self31;
reg [6:0] builder_sync_f_t_self32;
reg [7:0] builder_sync_f_t_self33;
reg [6:0] builder_sync_f_t_self34;
reg [7:0] builder_sync_f_t_self35;
reg [6:0] builder_sync_f_t_self36;
reg [7:0] builder_sync_f_t_self37;
reg [6:0] builder_sync_f_t_self38;
reg [7:0] builder_sync_f_t_self39;
reg [6:0] builder_sync_f_t_self40;
reg [7:0] builder_sync_f_t_self41;
reg [6:0] builder_sync_f_t_self42;
reg [7:0] builder_sync_f_t_self43;
reg [6:0] builder_sync_f_t_self44;
reg [7:0] builder_sync_f_t_self45;
reg [6:0] builder_sync_f_t_self46;
reg [7:0] builder_sync_f_t_self47;
reg [6:0] builder_sync_f_t_self48;
reg [7:0] builder_sync_f_t_self49;
reg [6:0] builder_sync_f_t_self50;
reg [7:0] builder_sync_f_t_self51;
reg [6:0] builder_sync_f_t_self52;
reg [7:0] builder_sync_f_t_self53;
reg [6:0] builder_sync_f_t_self54;
reg [7:0] builder_sync_f_t_self55;
reg [6:0] builder_sync_f_t_self56;
reg [7:0] builder_sync_f_t_self57;
reg [6:0] builder_sync_f_t_self58;
reg [31:0] builder_sync_rhs_self5;
reg [31:0] builder_sync_t_t_self0 = 32'd0;
reg [31:0] builder_sync_rhs_self6;
reg [31:0] builder_sync_t_t_self1 = 32'd0;
reg [31:0] builder_sync_t_rhs_self3;
reg builder_sync_t_rhs_self4;
reg builder_sync_t_rhs_self5;
reg builder_sync_t_rhs_self6;
reg builder_sync_t_rhs_self7;
reg builder_sync_t_rhs_self8;
reg builder_sync_t_rhs_self9;
reg builder_sync_t_rhs_self10;
reg builder_sync_t_rhs_self11;
reg builder_sync_t_rhs_self12;
reg builder_sync_t_rhs_self13;
reg builder_sync_t_rhs_self14;
reg builder_sync_t_rhs_self15;
reg builder_sync_t_rhs_self16;
reg builder_sync_t_rhs_self17;
reg builder_sync_t_rhs_self18;
reg builder_sync_t_rhs_self19;
reg [31:0] builder_sync_t_rhs_self20;
reg builder_sync_t_rhs_self21;
reg builder_sync_t_rhs_self22;
reg builder_sync_t_rhs_self23;
reg builder_sync_t_rhs_self24;
reg builder_sync_t_rhs_self25;
reg [31:0] builder_sync_t_rhs_self26;
reg builder_sync_t_rhs_self27;
reg builder_sync_t_rhs_self28;
reg builder_sync_t_rhs_self29;
reg builder_sync_t_rhs_self30;
reg builder_sync_t_rhs_self31;
reg builder_sync_t_rhs_self32;
reg builder_sync_t_rhs_self33;
reg builder_sync_t_rhs_self34;
reg [15:0] builder_sync_t_rhs_self35;
reg builder_sync_t_rhs_self36;
reg builder_sync_t_rhs_self37;
reg builder_sync_t_rhs_self38;
reg builder_sync_t_rhs_self39;
reg builder_sync_t_rhs_self40;
reg builder_sync_t_rhs_self41;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl00 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl01 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl10 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl11 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl0_async_reset;
wire builder_xilinxasyncresetsynchronizerimpl0_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl20 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl21 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl30 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl31 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl40 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl41 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl50 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl51 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl60 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl61 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl70 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl71 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl80 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl81 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl90 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl91 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl1_async_reset;
wire builder_xilinxasyncresetsynchronizerimpl1_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl2_async_reset;
wire builder_xilinxasyncresetsynchronizerimpl2_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl100 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl101 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl110 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl111 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl120 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl121 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl130 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl131 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl140 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl141 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl150 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl151 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl160 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl161 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl170 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl171 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl180 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl181 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl190 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl191 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl200 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl201 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl210 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl211 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl220 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl221 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl230 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl231 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl240 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl241 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl250 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl251 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl260 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl261 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl270 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl271 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl280 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl281 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl290 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl291 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl300 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl301 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl310 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl311 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl320 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl321 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl330 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl331 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl340 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl341 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl350 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl351 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl360 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl361 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl370 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl371 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl380 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl381 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl390 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl391 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl400 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl401 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl410 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl411 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl420 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl421 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl430 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl431 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl440 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl441 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl450 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl451 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl460 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl461 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl470 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl471 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl480 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl481 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl490 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl491 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl500 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl501 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl510 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl511 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl520 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl521 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl530 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl531 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl540 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl541 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl550 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl551 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl560 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl561 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl570 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl571 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl580 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl581 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl590 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl591 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl600 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl601 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl610 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl611 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl620 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl621 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl630 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl631 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl640 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl641 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl650 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl651 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl660 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl661 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl670 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl671 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl680 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl681 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl690 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl691 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl700 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl701 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl710 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl711 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl720 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl721 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl730 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl731 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl740 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl741 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl750 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl751 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl760 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl761 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl770 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl771 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl780 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl781 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl790 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl791 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl800 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl801 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl810 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl811 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl820 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl821 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl830 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl831 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl840 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl841 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl850 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl851 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl860 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl861 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl870 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl871 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl880 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl881 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl890 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl891 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl900 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl901 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl910 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl911 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl920 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl921 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl930 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl931 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl940 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl941 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl950 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl951 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl960 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl961 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl970 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl971 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl980 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl981 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl990 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl991 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1000 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1001 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1010 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1011 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1020 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1021 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1030 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1031 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1040 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1041 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1050 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1051 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1060 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1061 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1070 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1071 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1080 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1081 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1090 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1091 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1100 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1101 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1110 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1111 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1120 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1121 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1130 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1131 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1140 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1141 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1150 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1151 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1160 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1161 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1170 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1171 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1180 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1181 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1190 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1191 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1200 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1201 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1210 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1211 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1220 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1221 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1230 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1231 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1240 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1241 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1250 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1251 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1260 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1261 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1270 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1271 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1280 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1281 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1290 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1291 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1300 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1301 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1310 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1311 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1320 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1321 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1330 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1331 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1340 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1341 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1350 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1351 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1360 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1361 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1370 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1371 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1380 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1381 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1390 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1391 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1400 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1401 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1410 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1411 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1420 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1421 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1430 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1431 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1440 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1441 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1450 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1451 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1460 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1461 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1470 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1471 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1480 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1481 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1490 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1491 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1500 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1501 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1510 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1511 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1520 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1521 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1530 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1531 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1540 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1541 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1550 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1551 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1560 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1561 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1570 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1571 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1580 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1581 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1590 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1591 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1600 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1601 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1610 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1611 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1620 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1621 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1630 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1631 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1640 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1641 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1650 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1651 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1660 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1661 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1670 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1671 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1680 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1681 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1690 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1691 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1700 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1701 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1710 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1711 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1720 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1721 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1730 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1731 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1740 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1741 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1750 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1751 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1760 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1761 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1770 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1771 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1780 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl1781 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1790 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1791 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1800 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1801 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1810 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1811 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1820 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1821 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1830 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1831 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1840 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1841 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1850 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1851 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1860 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1861 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1870 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1871 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1880 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1881 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1890 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1891 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1900 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1901 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1910 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1911 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1920 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1921 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1930 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1931 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1940 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1941 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1950 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1951 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1960 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1961 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1970 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1971 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1980 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1981 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1990 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1991 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2000 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2001 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2010 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2011 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2020 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2021 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2030 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2031 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2040 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2041 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2050 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2051 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2060 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2061 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2070 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2071 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2080 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2081 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2090 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2091 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2100 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2101 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2110 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2111 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2120 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2121 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2130 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2131 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2140 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2141 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2150 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2151 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2160 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2161 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2170 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2171 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2180 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2181 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2190 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2191 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2200 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2201 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2210 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2211 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2220 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2221 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2230 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2231 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2240 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2241 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2250 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2251 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2260 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2261 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2270 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2271 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2280 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2281 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2290 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2291 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2300 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2301 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2310 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2311 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2320 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2321 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2330 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2331 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2340 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2341 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2350 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2351 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2360 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2361 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2370 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2371 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2380 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2381 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2390 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2391 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2400 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2401 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2410 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2411 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2420 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2421 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2430 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2431 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2440 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2441 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2450 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2451 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2460 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2461 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2470 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2471 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2480 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2481 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2490 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2491 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2500 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2501 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2510 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2511 = 1'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address = main_genericstandalone_genericstandalone_genericstandalone_master_p0_address;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank = main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cas_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cs_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_ras_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_we_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cke = main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_odt = main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_reset_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata = main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata = main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_valid = main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_valid;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address = main_genericstandalone_genericstandalone_genericstandalone_master_p1_address;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank = main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cas_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cs_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_ras_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_we_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cke = main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_odt = main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_reset_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata = main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata = main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_valid = main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_valid;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address = main_genericstandalone_genericstandalone_genericstandalone_master_p2_address;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank = main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cas_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cs_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_ras_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_we_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cke = main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_odt = main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_reset_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata = main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata = main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_valid = main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_valid;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address = main_genericstandalone_genericstandalone_genericstandalone_master_p3_address;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank = main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cas_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cs_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_ras_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_we_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cke = main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_odt = main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_reset_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata = main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata = main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_valid = main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_valid;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_address = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_bank;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cas_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cs_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cs_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_ras_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_we_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cke = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cke;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_odt = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_odt;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_reset_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_reset_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_mask;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata = main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata_valid = main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_valid;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_address = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_bank;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cas_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cs_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cs_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_ras_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_we_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cke = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cke;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_odt = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_odt;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_reset_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_reset_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_mask;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata = main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid = main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_valid;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_address = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_bank;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cas_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cs_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cs_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_ras_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_we_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cke = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cke;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_odt = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_odt;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_reset_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_reset_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_mask;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata = main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata_valid = main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_valid;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_address = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_bank;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cas_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cas_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cs_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cs_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_ras_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_ras_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_we_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_we_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cke = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cke;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_odt = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_odt;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_reset_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_reset_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_mask;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata = main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata_valid = main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_valid;
assign main_genericstandalone_virtual_led = main_genericstandalone_pcs_link_up;

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_interrupt <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_interrupt[0] <= main_genericstandalone_genericstandalone_genericstandalone_uart_irq;
	main_genericstandalone_genericstandalone_genericstandalone_interrupt[1] <= main_genericstandalone_genericstandalone_genericstandalone_timer0_irq;
	main_genericstandalone_genericstandalone_genericstandalone_interrupt[2] <= main_genericstandalone_sram166_irq;
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sram_we <= 8'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[0] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[0]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[1] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[1]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[2] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[2]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[3] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[3]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[4] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[4]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[5] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[5]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[6] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[6]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[7] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[7]);
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sram_adr = main_genericstandalone_genericstandalone_genericstandalone_sram_bus_adr[9:0];
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_sram_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w = main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_re;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_r;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_txfull_status = (~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_ack);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_last = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_last;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger = (~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_ack);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_ack;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_last = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_last;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rxempty_status = (~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_stb);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_w = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger = (~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_stb);

// synthesis translate_off
reg dummy_d_2;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_tx_clear <= 1'd0;
	if ((main_genericstandalone_genericstandalone_genericstandalone_uart_pending_re & main_genericstandalone_genericstandalone_genericstandalone_uart_pending_r[0])) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_2 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_3;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_status_w <= 2'd0;
	main_genericstandalone_genericstandalone_genericstandalone_uart_status_w[0] <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_status;
	main_genericstandalone_genericstandalone_genericstandalone_uart_status_w[1] <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_status;
// synthesis translate_off
	dummy_d_3 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_4;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear <= 1'd0;
	if ((main_genericstandalone_genericstandalone_genericstandalone_uart_pending_re & main_genericstandalone_genericstandalone_genericstandalone_uart_pending_r[1])) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_4 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_5;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w <= 2'd0;
	main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w[0] <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending;
	main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w[1] <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending;
// synthesis translate_off
	dummy_d_5 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_uart_irq = ((main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w[0] & main_genericstandalone_genericstandalone_genericstandalone_uart_storage[0]) | (main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w[1] & main_genericstandalone_genericstandalone_genericstandalone_uart_storage[1]));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_status = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_status = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_din = {main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_eop, main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_payload_data};
assign {main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_eop, main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_payload_data} = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_dout;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_readable;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_re = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_ack;

// synthesis translate_off
reg dummy_d_6;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr <= 4'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce - 1'd1);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_6 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_w = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_din;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_we = (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we & (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable | main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read = (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_readable & main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_re);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_adr = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_dout = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable = (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level != 5'd16);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_readable = (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level != 1'd0);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_din = {main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_eop, main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_payload_data};
assign {main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_eop, main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_payload_data} = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_dout;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_readable;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_re = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_ack;

// synthesis translate_off
reg dummy_d_7;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr <= 4'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce - 1'd1);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_7 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_w = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_din;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_we = (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we & (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable | main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read = (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_readable & main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_re);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_adr = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_dout = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable = (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level != 5'd16);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_readable = (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level != 1'd0);
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger = (main_genericstandalone_genericstandalone_genericstandalone_timer0_value != 1'd0);
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_status;

// synthesis translate_off
reg dummy_d_8;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_clear <= 1'd0;
	if ((main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_re & main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_r)) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_8 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending;
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_irq = (main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_w & main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage);
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_status = main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger;
assign main_genericstandalone_genericstandalone_crg_i_clk_sw = main_genericstandalone_rtiosyscrg_storage;

// synthesis translate_off
reg dummy_d_9;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_crg_reset <= 1'd0;
	builder_rtiosyscrg_next_state <= 2'd0;
	main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value0 <= 16'd0;
	main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value_ce0 <= 1'd0;
	main_genericstandalone_genericstandalone_crg_o_switch_rtiosyscrg_next_value1 <= 1'd0;
	main_genericstandalone_genericstandalone_crg_o_switch_rtiosyscrg_next_value_ce1 <= 1'd0;
	builder_rtiosyscrg_next_state <= builder_rtiosyscrg_state;
	case (builder_rtiosyscrg_state)
		1'd1: begin
			main_genericstandalone_genericstandalone_crg_reset <= 1'd1;
			if ((main_genericstandalone_genericstandalone_crg_delay_counter == 1'd0)) begin
				main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value0 <= 16'd65535;
				main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value_ce0 <= 1'd1;
				builder_rtiosyscrg_next_state <= 2'd2;
			end else begin
				main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value0 <= (main_genericstandalone_genericstandalone_crg_delay_counter - 1'd1);
				main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value_ce0 <= 1'd1;
			end
		end
		2'd2: begin
			main_genericstandalone_genericstandalone_crg_reset <= 1'd1;
			main_genericstandalone_genericstandalone_crg_o_switch_rtiosyscrg_next_value1 <= 1'd1;
			main_genericstandalone_genericstandalone_crg_o_switch_rtiosyscrg_next_value_ce1 <= 1'd1;
			main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value0 <= (main_genericstandalone_genericstandalone_crg_delay_counter - 1'd1);
			main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value_ce0 <= 1'd1;
			if ((main_genericstandalone_genericstandalone_crg_delay_counter == 1'd0)) begin
				builder_rtiosyscrg_next_state <= 1'd0;
			end
		end
		default: begin
			if ((main_genericstandalone_genericstandalone_crg_i_switch & (~main_genericstandalone_genericstandalone_crg_o_switch))) begin
				builder_rtiosyscrg_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_9 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtiosyscrg_async_reset = (((~main_genericstandalone_genericstandalone_crg_pll_locked) | (~main_genericstandalone_rtiosyscrg_mmcm_locked)) | main_genericstandalone_genericstandalone_crg_o_reset);
assign main_genericstandalone_genericstandalone_ddrphy_oe = ((main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en[1] | main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en[2]) | main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en[3]);

// synthesis translate_off
reg dummy_d_10;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_address <= 15'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_address <= 15'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_address <= 15'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_address <= 15'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en <= 1'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_storage[0]) begin
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_address <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_address <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_address <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_address <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_valid;
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_address <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_address <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_address <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_address <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_valid;
	end
// synthesis translate_off
	dummy_d_10 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cke = main_genericstandalone_genericstandalone_genericstandalone_storage[1];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cke = main_genericstandalone_genericstandalone_genericstandalone_storage[1];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cke = main_genericstandalone_genericstandalone_genericstandalone_storage[1];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cke = main_genericstandalone_genericstandalone_genericstandalone_storage[1];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_odt = main_genericstandalone_genericstandalone_genericstandalone_storage[2];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_odt = main_genericstandalone_genericstandalone_genericstandalone_storage[2];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_odt = main_genericstandalone_genericstandalone_genericstandalone_storage[2];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_odt = main_genericstandalone_genericstandalone_genericstandalone_storage[2];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_reset_n = main_genericstandalone_genericstandalone_genericstandalone_storage[3];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_reset_n = main_genericstandalone_genericstandalone_genericstandalone_storage[3];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_reset_n = main_genericstandalone_genericstandalone_genericstandalone_storage[3];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_reset_n = main_genericstandalone_genericstandalone_genericstandalone_storage[3];

// synthesis translate_off
reg dummy_d_11;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n <= 1'd1;
	if (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[0]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[1]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[2]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[3]);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_11 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_address = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_bank = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[4]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[5]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_12;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n <= 1'd1;
	if (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[0]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[1]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[2]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[3]);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_12 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_address = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_bank = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[4]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[5]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_13;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n <= 1'd1;
	if (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[0]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[1]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[2]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[3]);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_13 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_address = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_bank = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[4]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[5]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_14;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n <= 1'd1;
	if (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[0]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[1]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[2]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[3]);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_14 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_address = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_bank = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[4]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[5]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_mask = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset1 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset2 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset3 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset4 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset5 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset6 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset7 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];

// synthesis translate_off
reg dummy_d_15;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7 <= 1'd0;
	case (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7])
		1'd0: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0 <= 1'd1;
		end
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1 <= 1'd1;
		end
		2'd2: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2 <= 1'd1;
		end
		2'd3: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3 <= 1'd1;
		end
		3'd4: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4 <= 1'd1;
		end
		3'd5: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5 <= 1'd1;
		end
		3'd6: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6 <= 1'd1;
		end
		3'd7: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_15 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_hit = ((((((((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_idle = ((((((((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_wait = (~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write);
assign {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_swap_bank, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col_inc_next} = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col + 4'd8);
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read_ended = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_rdvalid_r & (~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_reset_n = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_odt = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cke = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cs_n = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_16;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address <= 15'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address <= 11'd1024;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
		end else begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read)) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col;
			end
		end
	end
// synthesis translate_off
	dummy_d_16 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_reset_n = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_odt = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cke = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cs_n = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_17;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address <= 15'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address <= 11'd1024;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
		end else begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read)) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col;
			end
		end
	end
// synthesis translate_off
	dummy_d_17 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_reset_n = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_odt = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cke = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cs_n = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_18;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address <= 15'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address <= 11'd1024;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
		end else begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read)) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col;
			end
		end
	end
// synthesis translate_off
	dummy_d_18 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_reset_n = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_odt = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cke = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cs_n = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_19;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address <= 15'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address <= 11'd1024;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
		end else begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read)) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col;
			end
		end
	end
// synthesis translate_off
	dummy_d_19 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r = {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata};
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_dat_w1 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_sel1 = (~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_sel);
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_done = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_count == 1'd0);

// synthesis translate_off
reg dummy_d_20;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_adr_inc <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_burst <= 1'd0;
	builder_minicon_next_state <= 6'd0;
	builder_minicon_next_state <= builder_minicon_state;
	case (builder_minicon_state)
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en <= 1'd1;
			builder_minicon_next_state <= 2'd2;
		end
		2'd2: begin
			if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= 1'd1;
				builder_minicon_next_state <= 1'd0;
			end
		end
		2'd3: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid;
			if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read_ended) begin
				builder_minicon_next_state <= 1'd0;
			end else begin
				if (((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti == 3'd7) & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack)) begin
					builder_minicon_next_state <= 3'd5;
				end
			end
		end
		3'd4: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_burst <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_adr_inc <= 1'd1;
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti == 3'd7)) begin
				builder_minicon_next_state <= 3'd5;
			end else begin
				if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_swap_bank) begin
					builder_minicon_next_state <= 2'd3;
				end
			end
		end
		3'd5: begin
			if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read_ended) begin
				builder_minicon_next_state <= 1'd0;
			end
		end
		3'd6: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= 1'd1;
			builder_minicon_next_state <= 4'd12;
		end
		3'd7: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_burst <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_adr_inc <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= 1'd1;
			if (((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti == 3'd7) | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_swap_bank)) begin
				builder_minicon_next_state <= 4'd12;
			end
		end
		4'd8: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd0;
			builder_minicon_next_state <= 5'd18;
		end
		4'd9: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n <= 1'd0;
			builder_minicon_next_state <= 4'd14;
		end
		4'd10: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n <= 1'd1;
			builder_minicon_next_state <= 5'd16;
		end
		4'd11: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd1;
			builder_minicon_next_state <= 5'd20;
		end
		4'd12: begin
			builder_minicon_next_state <= 4'd13;
		end
		4'd13: begin
			builder_minicon_next_state <= 1'd0;
		end
		4'd14: begin
			builder_minicon_next_state <= 4'd15;
		end
		4'd15: begin
			builder_minicon_next_state <= 4'd10;
		end
		5'd16: begin
			builder_minicon_next_state <= 5'd17;
		end
		5'd17: begin
			builder_minicon_next_state <= 1'd0;
		end
		5'd18: begin
			builder_minicon_next_state <= 5'd19;
		end
		5'd19: begin
			builder_minicon_next_state <= 4'd11;
		end
		5'd20: begin
			builder_minicon_next_state <= 5'd21;
		end
		5'd21: begin
			builder_minicon_next_state <= 5'd22;
		end
		5'd22: begin
			builder_minicon_next_state <= 5'd23;
		end
		5'd23: begin
			builder_minicon_next_state <= 5'd24;
		end
		5'd24: begin
			builder_minicon_next_state <= 5'd25;
		end
		5'd25: begin
			builder_minicon_next_state <= 5'd26;
		end
		5'd26: begin
			builder_minicon_next_state <= 5'd27;
		end
		5'd27: begin
			builder_minicon_next_state <= 5'd28;
		end
		5'd28: begin
			builder_minicon_next_state <= 5'd29;
		end
		5'd29: begin
			builder_minicon_next_state <= 5'd30;
		end
		5'd30: begin
			builder_minicon_next_state <= 5'd31;
		end
		5'd31: begin
			builder_minicon_next_state <= 6'd32;
		end
		6'd32: begin
			builder_minicon_next_state <= 6'd33;
		end
		6'd33: begin
			builder_minicon_next_state <= 6'd34;
		end
		6'd34: begin
			builder_minicon_next_state <= 6'd35;
		end
		6'd35: begin
			builder_minicon_next_state <= 6'd36;
		end
		6'd36: begin
			builder_minicon_next_state <= 6'd37;
		end
		6'd37: begin
			builder_minicon_next_state <= 6'd38;
		end
		6'd38: begin
			builder_minicon_next_state <= 6'd39;
		end
		6'd39: begin
			builder_minicon_next_state <= 6'd40;
		end
		6'd40: begin
			builder_minicon_next_state <= 6'd41;
		end
		6'd41: begin
			builder_minicon_next_state <= 6'd42;
		end
		6'd42: begin
			builder_minicon_next_state <= 6'd43;
		end
		6'd43: begin
			builder_minicon_next_state <= 6'd44;
		end
		6'd44: begin
			builder_minicon_next_state <= 6'd45;
		end
		6'd45: begin
			builder_minicon_next_state <= 6'd46;
		end
		6'd46: begin
			builder_minicon_next_state <= 6'd47;
		end
		6'd47: begin
			builder_minicon_next_state <= 6'd48;
		end
		6'd48: begin
			builder_minicon_next_state <= 6'd49;
		end
		6'd49: begin
			builder_minicon_next_state <= 6'd50;
		end
		6'd50: begin
			builder_minicon_next_state <= 6'd51;
		end
		6'd51: begin
			builder_minicon_next_state <= 6'd52;
		end
		6'd52: begin
			builder_minicon_next_state <= 1'd0;
		end
		default: begin
			if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_pending_refresh) begin
				builder_minicon_next_state <= 4'd8;
			end else begin
				if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_stb & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cyc)) begin
					if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_hit) begin
						if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_we) begin
							if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti == 2'd2)) begin
								builder_minicon_next_state <= 3'd7;
							end else begin
								builder_minicon_next_state <= 3'd6;
							end
						end else begin
							if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti == 2'd2)) begin
								builder_minicon_next_state <= 3'd4;
							end else begin
								builder_minicon_next_state <= 1'd1;
							end
						end
					end else begin
						if ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_idle)) begin
							if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_done) begin
								builder_minicon_next_state <= 4'd9;
							end
						end else begin
							builder_minicon_next_state <= 4'd10;
						end
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_20 <= dummy_s;
// synthesis translate_on
end
assign {main_genericstandalone_genericstandalone_genericstandalone_cache_newline, main_genericstandalone_genericstandalone_genericstandalone_cache_next_adr_offset} = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] + 1'd1);
assign main_genericstandalone_genericstandalone_genericstandalone_cache_last = (main_genericstandalone_genericstandalone_genericstandalone_cache_newline | (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cti != 2'd2));
assign main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_adr = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[13:3];

// synthesis translate_off
reg dummy_d_21;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_we <= 64'd0;
	main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_w <= 512'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_cache_write_from_slave) begin
		main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_w <= {4{main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_r}};
		main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_we <= {({16{(main_genericstandalone_genericstandalone_genericstandalone_cache == 1'd0)}} & {16{1'd1}}), ({16{(main_genericstandalone_genericstandalone_genericstandalone_cache == 1'd1)}} & {16{1'd1}}), ({16{(main_genericstandalone_genericstandalone_genericstandalone_cache == 2'd2)}} & {16{1'd1}}), ({16{(main_genericstandalone_genericstandalone_genericstandalone_cache == 2'd3)}} & {16{1'd1}})};
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_w <= {8{main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_w}};
		if ((((main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cyc & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_stb) & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_we) & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack)) begin
			main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_we <= {({8{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] == 1'd0)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({8{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] == 1'd1)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({8{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] == 2'd2)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({8{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] == 2'd3)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({8{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] == 3'd4)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({8{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] == 3'd5)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({8{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] == 3'd6)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({8{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0] == 3'd7)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel)};
		end
	end
// synthesis translate_off
	dummy_d_21 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_22;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w <= 128'd0;
	case (main_genericstandalone_genericstandalone_genericstandalone_cache)
		1'd0: begin
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[511:384];
		end
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[383:256];
		end
		2'd2: begin
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[255:128];
		end
		default: begin
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[127:0];
		end
	endcase
// synthesis translate_off
	dummy_d_22 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_sel = 16'd65535;

// synthesis translate_off
reg dummy_d_23;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= 64'd0;
	case (main_genericstandalone_genericstandalone_genericstandalone_cache_adr_offset_r)
		1'd0: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[511:448];
		end
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[447:384];
		end
		2'd2: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[383:320];
		end
		2'd3: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[319:256];
		end
		3'd4: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[255:192];
		end
		3'd5: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[191:128];
		end
		3'd6: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[127:64];
		end
		default: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r[63:0];
		end
	endcase
// synthesis translate_off
	dummy_d_23 <= dummy_s;
// synthesis translate_on
end
assign {main_genericstandalone_genericstandalone_genericstandalone_cache_tag_do_dirty, main_genericstandalone_genericstandalone_genericstandalone_cache_tag_do_tag} = main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_dat_w = {main_genericstandalone_genericstandalone_genericstandalone_cache_tag_di_dirty, main_genericstandalone_genericstandalone_genericstandalone_cache_tag_di_tag};
assign main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_adr = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[13:3];
assign main_genericstandalone_genericstandalone_genericstandalone_cache_tag_di_tag = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[28:14];
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_adr = {main_genericstandalone_genericstandalone_genericstandalone_cache_tag_do_tag, main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[13:3], main_genericstandalone_genericstandalone_genericstandalone_cache};

// synthesis translate_off
reg dummy_d_24;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cti <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_cache_write_from_slave <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_cache_adr_inc <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_we <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_cache_tag_di_dirty <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_cache_word_clr <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_cache_word_inc <= 1'd0;
	builder_cache_next_state <= 3'd0;
	builder_cache_next_state <= builder_cache_state;
	case (builder_cache_state)
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_cache_word_clr <= 1'd1;
			if ((main_genericstandalone_genericstandalone_genericstandalone_cache_tag_do_tag == main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[28:14])) begin
				main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack <= 1'd1;
				main_genericstandalone_genericstandalone_genericstandalone_cache_adr_inc <= 1'd1;
				if (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_we) begin
					main_genericstandalone_genericstandalone_genericstandalone_cache_tag_di_dirty <= 1'd1;
					main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_we <= 1'd1;
				end
				if (main_genericstandalone_genericstandalone_genericstandalone_cache_last) begin
					builder_cache_next_state <= 1'd0;
				end
			end else begin
				if (main_genericstandalone_genericstandalone_genericstandalone_cache_tag_do_dirty) begin
					builder_cache_next_state <= 2'd2;
				end else begin
					builder_cache_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cti <= ((main_genericstandalone_genericstandalone_genericstandalone_cache == 2'd3) ? 3'd7 : 2'd2);
			if (main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack) begin
				main_genericstandalone_genericstandalone_genericstandalone_cache_word_inc <= 1'd1;
				if ((main_genericstandalone_genericstandalone_genericstandalone_cache == 2'd3)) begin
					builder_cache_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_we <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_cache_word_clr <= 1'd1;
			builder_cache_next_state <= 3'd4;
		end
		3'd4: begin
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cti <= ((main_genericstandalone_genericstandalone_genericstandalone_cache == 2'd3) ? 3'd7 : 2'd2);
			if (main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack) begin
				main_genericstandalone_genericstandalone_genericstandalone_cache_write_from_slave <= 1'd1;
				main_genericstandalone_genericstandalone_genericstandalone_cache_word_inc <= 1'd1;
				if ((main_genericstandalone_genericstandalone_genericstandalone_cache == 2'd3)) begin
					builder_cache_next_state <= 1'd1;
				end else begin
					builder_cache_next_state <= 3'd4;
				end
			end
		end
		default: begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cyc & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_stb)) begin
				builder_cache_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_24 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_virtual_leds_status[0] = main_genericstandalone_virtual_led;
assign main_genericstandalone_genericstandalone_spiflash_bus_dat_r = {main_genericstandalone_genericstandalone_spiflash_sr[7:0], main_genericstandalone_genericstandalone_spiflash_sr[15:8], main_genericstandalone_genericstandalone_spiflash_sr[23:16], main_genericstandalone_genericstandalone_spiflash_sr[31:24], main_genericstandalone_genericstandalone_spiflash_sr[39:32], main_genericstandalone_genericstandalone_spiflash_sr[47:40], main_genericstandalone_genericstandalone_spiflash_sr[55:48], main_genericstandalone_genericstandalone_spiflash_sr[63:56]};

// synthesis translate_off
reg dummy_d_25;
// synthesis translate_on
always @(*) begin
	spiflash2x_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_clk <= 1'd0;
	main_genericstandalone_genericstandalone_spiflash_status <= 1'd0;
	main_genericstandalone_genericstandalone_spiflash_o <= 2'd0;
	main_genericstandalone_genericstandalone_spiflash_oe <= 1'd0;
	if (main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage) begin
		main_genericstandalone_genericstandalone_clk <= main_genericstandalone_genericstandalone_spiflash_bitbang_storage[1];
		spiflash2x_cs_n <= main_genericstandalone_genericstandalone_spiflash_bitbang_storage[2];
		if (main_genericstandalone_genericstandalone_spiflash_bitbang_storage[3]) begin
			main_genericstandalone_genericstandalone_spiflash_oe <= 1'd0;
		end else begin
			main_genericstandalone_genericstandalone_spiflash_oe <= 1'd1;
		end
		if (main_genericstandalone_genericstandalone_spiflash_bitbang_storage[1]) begin
			main_genericstandalone_genericstandalone_spiflash_status <= main_genericstandalone_genericstandalone_spiflash_i0[1];
		end
		main_genericstandalone_genericstandalone_spiflash_o <= {{1{1'd1}}, main_genericstandalone_genericstandalone_spiflash_bitbang_storage[0]};
	end else begin
		main_genericstandalone_genericstandalone_clk <= main_genericstandalone_genericstandalone_spiflash_clk;
		spiflash2x_cs_n <= main_genericstandalone_genericstandalone_spiflash_cs_n;
		main_genericstandalone_genericstandalone_spiflash_o <= main_genericstandalone_genericstandalone_spiflash_sr[63:62];
		main_genericstandalone_genericstandalone_spiflash_oe <= main_genericstandalone_genericstandalone_spiflash_dq_oe;
	end
// synthesis translate_off
	dummy_d_25 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_icap_counter_rst = (main_genericstandalone_genericstandalone_icap_counter0 == 1'd0);
assign main_genericstandalone_genericstandalone_icap_i = main_genericstandalone_genericstandalone_icap_iprog_re;
assign main_genericstandalone_genericstandalone_icap_o = (main_genericstandalone_genericstandalone_icap_toggle_o ^ main_genericstandalone_genericstandalone_icap_toggle_o_r);

// synthesis translate_off
reg dummy_d_26;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_icap_icap_csib <= 1'd0;
	main_genericstandalone_genericstandalone_icap_icap_i <= 32'd0;
	main_genericstandalone_genericstandalone_icap_icap_rdwrb <= 1'd0;
	builder_icap_next_state <= 1'd0;
	main_genericstandalone_genericstandalone_icap_counter1_icap_next_value <= 4'd0;
	main_genericstandalone_genericstandalone_icap_counter1_icap_next_value_ce <= 1'd0;
	builder_icap_next_state <= builder_icap_state;
	case (builder_icap_state)
		1'd1: begin
			main_genericstandalone_genericstandalone_icap_icap_rdwrb <= 1'd0;
			main_genericstandalone_genericstandalone_icap_icap_csib <= 1'd0;
			main_genericstandalone_genericstandalone_icap_icap_i <= builder_comb_basiclowerer_self;
			main_genericstandalone_genericstandalone_icap_counter1_icap_next_value <= (main_genericstandalone_genericstandalone_icap_counter1 + 1'd1);
			main_genericstandalone_genericstandalone_icap_counter1_icap_next_value_ce <= 1'd1;
			if ((main_genericstandalone_genericstandalone_icap_counter1 == 4'd10)) begin
				builder_icap_next_state <= 1'd0;
			end else begin
				builder_icap_next_state <= 1'd1;
			end
		end
		default: begin
			main_genericstandalone_genericstandalone_icap_icap_rdwrb <= 1'd1;
			main_genericstandalone_genericstandalone_icap_icap_csib <= 1'd1;
			if (main_genericstandalone_genericstandalone_icap_o) begin
				builder_icap_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_26 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_qpll_reset = main_genericstandalone_tx_init_qpll_reset0;
assign main_genericstandalone_tx_init_qpll_lock0 = main_genericstandalone_genericstandalone_qpll_lock;
assign main_genericstandalone_tx_reset = main_genericstandalone_tx_init_tx_reset0;
assign main_genericstandalone_rx_init_enable = main_genericstandalone_tx_init_done;
assign main_genericstandalone_rx_reset = main_genericstandalone_rx_init_rx_reset0;
assign main_genericstandalone_rx_init_rx_pma_reset_done0 = main_genericstandalone_rx_pma_reset_done;
assign main_genericstandalone_drpaddr = main_genericstandalone_rx_init_drpaddr;
assign main_genericstandalone_drpen = main_genericstandalone_rx_init_drpen;
assign main_genericstandalone_drpdi = main_genericstandalone_rx_init_drpdi;
assign main_genericstandalone_rx_init_drprdy = main_genericstandalone_drprdy;
assign main_genericstandalone_rx_init_drpdo = main_genericstandalone_drpdo;
assign main_genericstandalone_drpwe = main_genericstandalone_rx_init_drpwe;
assign main_genericstandalone_i = main_genericstandalone_pcs_restart;
assign main_genericstandalone_rx_init_restart = main_genericstandalone_o;
assign main_genericstandalone_tx_data0 = main_genericstandalone_tx_data_half;
assign main_genericstandalone_rx_data_half = main_genericstandalone_rx_data0;
assign main_genericstandalone_tx_data1 = main_genericstandalone_pcs_transmitpath_encoder2;
assign main_genericstandalone_pcs_receivepath_input = main_genericstandalone_rx_data1;
assign main_genericstandalone_pcs_transmitpath_tx_stb = main_genericstandalone_pcs_sink_stb;
assign main_genericstandalone_pcs_sink_ack = main_genericstandalone_pcs_transmitpath_tx_ack;
assign main_genericstandalone_pcs_transmitpath_tx_data = main_genericstandalone_pcs_sink_payload_data;
assign main_genericstandalone_pcs_source_eop = ((~main_genericstandalone_pcs_receivepath_rx_en) & main_genericstandalone_pcs_rx_en_d);
assign main_genericstandalone_pcs_seen_valid_ci_i = main_genericstandalone_pcs_receivepath_seen_valid_ci;
assign main_genericstandalone_pcs_is_sgmii = main_genericstandalone_pcs_lp_abi_o[0];
assign main_genericstandalone_pcs_linkdown = ((main_genericstandalone_pcs_lp_abi_o[0] & (~main_genericstandalone_pcs_lp_abi_o[15])) | (main_genericstandalone_pcs_lp_abi_o == 1'd0));
assign main_genericstandalone_pcs_transmitpath_sgmii_speed = (main_genericstandalone_pcs_lp_abi_o[0] ? main_genericstandalone_pcs_lp_abi_o[11:10] : 2'd2);
assign main_genericstandalone_pcs_receivepath_sgmii_speed = (main_genericstandalone_pcs_lp_abi_i[0] ? main_genericstandalone_pcs_lp_abi_i[11:10] : 2'd2);
assign main_genericstandalone_pcs_transmitpath_config_reg = (main_genericstandalone_pcs_tx_config_empty ? 1'd0 : (((((main_genericstandalone_pcs_is_sgmii | ((~main_genericstandalone_pcs_is_sgmii) <<< 3'd5)) | ((main_genericstandalone_pcs_lp_abi_o[0] ? main_genericstandalone_pcs_lp_abi_o[11:10] : 1'd0) <<< 4'd10)) | (main_genericstandalone_pcs_is_sgmii <<< 4'd12)) | (main_genericstandalone_pcs_autoneg_ack <<< 4'd14)) | (main_genericstandalone_pcs_is_sgmii & main_genericstandalone_pcs_link_up)));
assign main_genericstandalone_pcs_transmitpath_encoder_d = main_genericstandalone_pcs_transmitpath_encoder0;
assign main_genericstandalone_pcs_transmitpath_encoder_k = main_genericstandalone_pcs_transmitpath_encoder1;
assign main_genericstandalone_pcs_transmitpath_encoder_disp_inter = (main_genericstandalone_pcs_transmitpath_encoder_disp_in ^ main_genericstandalone_pcs_transmitpath_encoder_code6b_unbalanced);

// synthesis translate_off
reg dummy_d_27;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_encoder_output_6b <= 6'd0;
	if (((~main_genericstandalone_pcs_transmitpath_encoder_disp_in) & main_genericstandalone_pcs_transmitpath_encoder_code6b_flip)) begin
		main_genericstandalone_pcs_transmitpath_encoder_output_6b <= (~main_genericstandalone_pcs_transmitpath_encoder_code6b);
	end else begin
		main_genericstandalone_pcs_transmitpath_encoder_output_6b <= main_genericstandalone_pcs_transmitpath_encoder_code6b;
	end
// synthesis translate_off
	dummy_d_27 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_28;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_encoder_disp_out <= 1'd0;
	main_genericstandalone_pcs_transmitpath_encoder_output_4b <= 4'd0;
	if (((~main_genericstandalone_pcs_transmitpath_encoder_disp_inter) & main_genericstandalone_pcs_transmitpath_encoder_alt7_rd0)) begin
		main_genericstandalone_pcs_transmitpath_encoder_disp_out <= (~main_genericstandalone_pcs_transmitpath_encoder_disp_inter);
		main_genericstandalone_pcs_transmitpath_encoder_output_4b <= 3'd7;
	end else begin
		if ((main_genericstandalone_pcs_transmitpath_encoder_disp_inter & main_genericstandalone_pcs_transmitpath_encoder_alt7_rd1)) begin
			main_genericstandalone_pcs_transmitpath_encoder_disp_out <= (~main_genericstandalone_pcs_transmitpath_encoder_disp_inter);
			main_genericstandalone_pcs_transmitpath_encoder_output_4b <= 4'd8;
		end else begin
			main_genericstandalone_pcs_transmitpath_encoder_disp_out <= (main_genericstandalone_pcs_transmitpath_encoder_disp_inter ^ main_genericstandalone_pcs_transmitpath_encoder_code4b_unbalanced);
			if (((~main_genericstandalone_pcs_transmitpath_encoder_disp_inter) & main_genericstandalone_pcs_transmitpath_encoder_code4b_flip)) begin
				main_genericstandalone_pcs_transmitpath_encoder_output_4b <= (~main_genericstandalone_pcs_transmitpath_encoder_code4b);
			end else begin
				main_genericstandalone_pcs_transmitpath_encoder_output_4b <= main_genericstandalone_pcs_transmitpath_encoder_code4b;
			end
		end
	end
// synthesis translate_off
	dummy_d_28 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_pcs_transmitpath_encoder_output_msb_first = {main_genericstandalone_pcs_transmitpath_encoder_output_6b, main_genericstandalone_pcs_transmitpath_encoder_output_4b};

// synthesis translate_off
reg dummy_d_29;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_encoder_output <= 10'd0;
	main_genericstandalone_pcs_transmitpath_encoder_output[0] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[9];
	main_genericstandalone_pcs_transmitpath_encoder_output[1] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[8];
	main_genericstandalone_pcs_transmitpath_encoder_output[2] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[7];
	main_genericstandalone_pcs_transmitpath_encoder_output[3] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[6];
	main_genericstandalone_pcs_transmitpath_encoder_output[4] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[5];
	main_genericstandalone_pcs_transmitpath_encoder_output[5] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[4];
	main_genericstandalone_pcs_transmitpath_encoder_output[6] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[3];
	main_genericstandalone_pcs_transmitpath_encoder_output[7] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[2];
	main_genericstandalone_pcs_transmitpath_encoder_output[8] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[1];
	main_genericstandalone_pcs_transmitpath_encoder_output[9] <= main_genericstandalone_pcs_transmitpath_encoder_output_msb_first[0];
// synthesis translate_off
	dummy_d_29 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_30;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_tx_ack <= 1'd0;
	main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd0;
	main_genericstandalone_pcs_transmitpath_encoder1 <= 1'd0;
	main_genericstandalone_pcs_transmitpath_load_config_reg_buffer <= 1'd0;
	main_genericstandalone_pcs_transmitpath_timer_en <= 1'd0;
	builder_a7_1000basex_transmitpath_next_state <= 3'd0;
	main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value <= 1'd0;
	main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value_ce <= 1'd0;
	builder_a7_1000basex_transmitpath_next_state <= builder_a7_1000basex_transmitpath_state;
	case (builder_a7_1000basex_transmitpath_state)
		1'd1: begin
			if (main_genericstandalone_pcs_transmitpath_c_type) begin
				main_genericstandalone_pcs_transmitpath_encoder0 <= 7'd66;
			end else begin
				main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd181;
			end
			main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value <= (~main_genericstandalone_pcs_transmitpath_c_type);
			main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value_ce <= 1'd1;
			builder_a7_1000basex_transmitpath_next_state <= 2'd2;
		end
		2'd2: begin
			main_genericstandalone_pcs_transmitpath_encoder0 <= main_genericstandalone_pcs_transmitpath_config_reg_buffer[7:0];
			builder_a7_1000basex_transmitpath_next_state <= 2'd3;
		end
		2'd3: begin
			main_genericstandalone_pcs_transmitpath_encoder0 <= main_genericstandalone_pcs_transmitpath_config_reg_buffer[15:8];
			builder_a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		3'd4: begin
			if (main_genericstandalone_pcs_transmitpath_encoder3) begin
				main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd197;
			end else begin
				main_genericstandalone_pcs_transmitpath_encoder0 <= 7'd80;
			end
			builder_a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		3'd5: begin
			if (main_genericstandalone_pcs_transmitpath_tx_stb) begin
				main_genericstandalone_pcs_transmitpath_tx_ack <= (main_genericstandalone_pcs_transmitpath_timer == 1'd0);
				main_genericstandalone_pcs_transmitpath_timer_en <= 1'd1;
				main_genericstandalone_pcs_transmitpath_encoder0 <= main_genericstandalone_pcs_transmitpath_tx_data;
			end else begin
				main_genericstandalone_pcs_transmitpath_tx_ack <= 1'd1;
				main_genericstandalone_pcs_transmitpath_encoder1 <= 1'd1;
				main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd253;
				builder_a7_1000basex_transmitpath_next_state <= 3'd6;
			end
		end
		3'd6: begin
			main_genericstandalone_pcs_transmitpath_encoder1 <= 1'd1;
			main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd247;
			if (main_genericstandalone_pcs_transmitpath_parity) begin
				builder_a7_1000basex_transmitpath_next_state <= 1'd0;
			end else begin
				builder_a7_1000basex_transmitpath_next_state <= 3'd7;
			end
		end
		3'd7: begin
			main_genericstandalone_pcs_transmitpath_encoder1 <= 1'd1;
			main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd247;
			builder_a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		default: begin
			if (main_genericstandalone_pcs_transmitpath_config_stb) begin
				main_genericstandalone_pcs_transmitpath_tx_ack <= 1'd1;
				main_genericstandalone_pcs_transmitpath_load_config_reg_buffer <= 1'd1;
				main_genericstandalone_pcs_transmitpath_encoder1 <= 1'd1;
				main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd188;
				builder_a7_1000basex_transmitpath_next_state <= 1'd1;
			end else begin
				if (main_genericstandalone_pcs_transmitpath_tx_stb) begin
					main_genericstandalone_pcs_transmitpath_tx_ack <= (main_genericstandalone_pcs_transmitpath_timer == 1'd0);
					main_genericstandalone_pcs_transmitpath_timer_en <= 1'd1;
					main_genericstandalone_pcs_transmitpath_encoder1 <= 1'd1;
					main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd251;
					builder_a7_1000basex_transmitpath_next_state <= 3'd5;
				end else begin
					main_genericstandalone_pcs_transmitpath_tx_ack <= 1'd1;
					main_genericstandalone_pcs_transmitpath_encoder1 <= 1'd1;
					main_genericstandalone_pcs_transmitpath_encoder0 <= 8'd188;
					builder_a7_1000basex_transmitpath_next_state <= 3'd4;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_30 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_pcs_receivepath_rx_data = (main_genericstandalone_pcs_receivepath_first_preamble_byte ? 7'd85 : main_genericstandalone_pcs_receivepath_d);
assign main_genericstandalone_pcs_receivepath_sample_en = (main_genericstandalone_pcs_receivepath_rx_en & (main_genericstandalone_pcs_receivepath_timer == 1'd0));

// synthesis translate_off
reg dummy_d_31;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_receivepath_input_msb_first <= 10'd0;
	main_genericstandalone_pcs_receivepath_input_msb_first[0] <= main_genericstandalone_pcs_receivepath_input[9];
	main_genericstandalone_pcs_receivepath_input_msb_first[1] <= main_genericstandalone_pcs_receivepath_input[8];
	main_genericstandalone_pcs_receivepath_input_msb_first[2] <= main_genericstandalone_pcs_receivepath_input[7];
	main_genericstandalone_pcs_receivepath_input_msb_first[3] <= main_genericstandalone_pcs_receivepath_input[6];
	main_genericstandalone_pcs_receivepath_input_msb_first[4] <= main_genericstandalone_pcs_receivepath_input[5];
	main_genericstandalone_pcs_receivepath_input_msb_first[5] <= main_genericstandalone_pcs_receivepath_input[4];
	main_genericstandalone_pcs_receivepath_input_msb_first[6] <= main_genericstandalone_pcs_receivepath_input[3];
	main_genericstandalone_pcs_receivepath_input_msb_first[7] <= main_genericstandalone_pcs_receivepath_input[2];
	main_genericstandalone_pcs_receivepath_input_msb_first[8] <= main_genericstandalone_pcs_receivepath_input[1];
	main_genericstandalone_pcs_receivepath_input_msb_first[9] <= main_genericstandalone_pcs_receivepath_input[0];
// synthesis translate_off
	dummy_d_31 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_pcs_receivepath_d = {main_genericstandalone_pcs_receivepath_code3b, main_genericstandalone_pcs_receivepath_code5b};

// synthesis translate_off
reg dummy_d_32;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_receivepath_rx_en <= 1'd0;
	main_genericstandalone_pcs_receivepath_seen_valid_ci <= 1'd0;
	main_genericstandalone_pcs_receivepath_load_config_reg_lsb <= 1'd0;
	main_genericstandalone_pcs_receivepath_load_config_reg_msb <= 1'd0;
	main_genericstandalone_pcs_receivepath_first_preamble_byte <= 1'd0;
	main_genericstandalone_pcs_receivepath_timer_en <= 1'd0;
	builder_a7_1000basex_receivepath_next_state <= 3'd0;
	builder_a7_1000basex_receivepath_next_state <= builder_a7_1000basex_receivepath_state;
	case (builder_a7_1000basex_receivepath_state)
		1'd1: begin
			builder_a7_1000basex_receivepath_next_state <= 1'd0;
			if ((~main_genericstandalone_pcs_receivepath_k)) begin
				if (((main_genericstandalone_pcs_receivepath_d == 8'd181) | (main_genericstandalone_pcs_receivepath_d == 7'd66))) begin
					main_genericstandalone_pcs_receivepath_seen_valid_ci <= 1'd1;
					builder_a7_1000basex_receivepath_next_state <= 2'd2;
				end
				if (((main_genericstandalone_pcs_receivepath_d == 8'd197) | (main_genericstandalone_pcs_receivepath_d == 7'd80))) begin
					main_genericstandalone_pcs_receivepath_seen_valid_ci <= 1'd1;
					builder_a7_1000basex_receivepath_next_state <= 1'd0;
				end
			end
		end
		2'd2: begin
			if (main_genericstandalone_pcs_receivepath_k) begin
				if ((main_genericstandalone_pcs_receivepath_d == 8'd251)) begin
					main_genericstandalone_pcs_receivepath_rx_en <= 1'd1;
					main_genericstandalone_pcs_receivepath_timer_en <= 1'd1;
					main_genericstandalone_pcs_receivepath_first_preamble_byte <= 1'd1;
					builder_a7_1000basex_receivepath_next_state <= 3'd4;
				end else begin
					builder_a7_1000basex_receivepath_next_state <= 1'd0;
				end
			end else begin
				main_genericstandalone_pcs_receivepath_load_config_reg_lsb <= 1'd1;
				builder_a7_1000basex_receivepath_next_state <= 2'd3;
			end
		end
		2'd3: begin
			if ((~main_genericstandalone_pcs_receivepath_k)) begin
				main_genericstandalone_pcs_receivepath_load_config_reg_msb <= 1'd1;
			end
			builder_a7_1000basex_receivepath_next_state <= 1'd0;
		end
		3'd4: begin
			if (main_genericstandalone_pcs_receivepath_k) begin
				builder_a7_1000basex_receivepath_next_state <= 1'd0;
			end else begin
				main_genericstandalone_pcs_receivepath_rx_en <= 1'd1;
				main_genericstandalone_pcs_receivepath_timer_en <= 1'd1;
			end
		end
		default: begin
			if (main_genericstandalone_pcs_receivepath_k) begin
				if ((main_genericstandalone_pcs_receivepath_d == 8'd188)) begin
					builder_a7_1000basex_receivepath_next_state <= 1'd1;
				end
				if ((main_genericstandalone_pcs_receivepath_d == 8'd251)) begin
					main_genericstandalone_pcs_receivepath_rx_en <= 1'd1;
					main_genericstandalone_pcs_receivepath_timer_en <= 1'd1;
					main_genericstandalone_pcs_receivepath_first_preamble_byte <= 1'd1;
					builder_a7_1000basex_receivepath_next_state <= 3'd4;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_32 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_pcs_lp_abi_wait = (~main_genericstandalone_pcs_lp_abi_ping_i);
assign main_genericstandalone_pcs_lp_abi_ping_i = ((main_genericstandalone_pcs_lp_abi_starter | main_genericstandalone_pcs_lp_abi_pong_o) | main_genericstandalone_pcs_lp_abi_done);
assign main_genericstandalone_pcs_lp_abi_pong_i = main_genericstandalone_pcs_lp_abi_ping_o1;
assign main_genericstandalone_pcs_lp_abi_ping_o0 = (main_genericstandalone_pcs_lp_abi_ping_toggle_o ^ main_genericstandalone_pcs_lp_abi_ping_toggle_o_r);
assign main_genericstandalone_pcs_lp_abi_pong_o = (main_genericstandalone_pcs_lp_abi_pong_toggle_o ^ main_genericstandalone_pcs_lp_abi_pong_toggle_o_r);
assign main_genericstandalone_pcs_lp_abi_done = (main_genericstandalone_pcs_lp_abi_count == 1'd0);
assign main_genericstandalone_pcs_seen_valid_ci_o = (main_genericstandalone_pcs_seen_valid_ci_toggle_o ^ main_genericstandalone_pcs_seen_valid_ci_toggle_o_r);
assign main_genericstandalone_pcs_rx_config_reg_abi_o = (main_genericstandalone_pcs_rx_config_reg_abi_toggle_o ^ main_genericstandalone_pcs_rx_config_reg_abi_toggle_o_r);
assign main_genericstandalone_pcs_rx_config_reg_ack_o = (main_genericstandalone_pcs_rx_config_reg_ack_toggle_o ^ main_genericstandalone_pcs_rx_config_reg_ack_toggle_o_r);
assign main_genericstandalone_pcs_waittimer0_done = (main_genericstandalone_pcs_waittimer0_count == 1'd0);
assign main_genericstandalone_pcs_waittimer1_done = (main_genericstandalone_pcs_waittimer1_count == 1'd0);

// synthesis translate_off
reg dummy_d_33;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_config_stb <= 1'd0;
	main_genericstandalone_pcs_link_up <= 1'd0;
	main_genericstandalone_pcs_restart <= 1'd0;
	main_genericstandalone_pcs_tx_config_empty <= 1'd0;
	main_genericstandalone_pcs_autoneg_ack <= 1'd0;
	main_genericstandalone_pcs_waittimer0_wait <= 1'd0;
	main_genericstandalone_pcs_waittimer1_wait <= 1'd0;
	builder_a7_1000basex_fsm_next_state <= 3'd0;
	builder_a7_1000basex_fsm_next_state <= builder_a7_1000basex_fsm_state;
	case (builder_a7_1000basex_fsm_state)
		1'd1: begin
			main_genericstandalone_pcs_transmitpath_config_stb <= 1'd1;
			if (main_genericstandalone_pcs_rx_config_reg_abi_o) begin
				builder_a7_1000basex_fsm_next_state <= 2'd2;
			end
			if ((main_genericstandalone_pcs_checker_tick & (~main_genericstandalone_pcs_checker_ok))) begin
				main_genericstandalone_pcs_restart <= 1'd1;
				builder_a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		2'd2: begin
			main_genericstandalone_pcs_transmitpath_config_stb <= 1'd1;
			main_genericstandalone_pcs_autoneg_ack <= 1'd1;
			if (main_genericstandalone_pcs_rx_config_reg_ack_o) begin
				builder_a7_1000basex_fsm_next_state <= 2'd3;
			end
			if ((main_genericstandalone_pcs_checker_tick & (~main_genericstandalone_pcs_checker_ok))) begin
				main_genericstandalone_pcs_restart <= 1'd1;
				builder_a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		2'd3: begin
			main_genericstandalone_pcs_transmitpath_config_stb <= 1'd1;
			main_genericstandalone_pcs_autoneg_ack <= 1'd1;
			main_genericstandalone_pcs_waittimer0_wait <= (~main_genericstandalone_pcs_is_sgmii);
			main_genericstandalone_pcs_waittimer1_wait <= main_genericstandalone_pcs_is_sgmii;
			if (((main_genericstandalone_pcs_is_sgmii & main_genericstandalone_pcs_waittimer1_done) | ((~main_genericstandalone_pcs_is_sgmii) & main_genericstandalone_pcs_waittimer0_done))) begin
				builder_a7_1000basex_fsm_next_state <= 3'd4;
			end
			if ((main_genericstandalone_pcs_checker_tick & (~main_genericstandalone_pcs_checker_ok))) begin
				main_genericstandalone_pcs_restart <= 1'd1;
				builder_a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		3'd4: begin
			main_genericstandalone_pcs_link_up <= 1'd1;
			if (((main_genericstandalone_pcs_checker_tick & (~main_genericstandalone_pcs_checker_ok)) | main_genericstandalone_pcs_linkdown)) begin
				main_genericstandalone_pcs_restart <= 1'd1;
				builder_a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_pcs_transmitpath_config_stb <= 1'd1;
			main_genericstandalone_pcs_tx_config_empty <= 1'd1;
			main_genericstandalone_pcs_waittimer0_wait <= 1'd1;
			if (main_genericstandalone_pcs_waittimer0_done) begin
				builder_a7_1000basex_fsm_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_33 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_34;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_init_done <= 1'd0;
	main_genericstandalone_tx_init_qpll_reset1 <= 1'd0;
	main_genericstandalone_tx_init_tx_reset1 <= 1'd0;
	builder_a7_1000basex_gtptxinit_next_state <= 2'd0;
	builder_a7_1000basex_gtptxinit_next_state <= builder_a7_1000basex_gtptxinit_state;
	case (builder_a7_1000basex_gtptxinit_state)
		1'd1: begin
			main_genericstandalone_tx_init_tx_reset1 <= 1'd1;
			main_genericstandalone_tx_init_qpll_reset1 <= 1'd1;
			if (main_genericstandalone_tx_init_tick) begin
				builder_a7_1000basex_gtptxinit_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_genericstandalone_tx_init_tx_reset1 <= 1'd1;
			if ((main_genericstandalone_tx_init_qpll_lock1 & main_genericstandalone_tx_init_tick)) begin
				builder_a7_1000basex_gtptxinit_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_genericstandalone_tx_init_done <= 1'd1;
		end
		default: begin
			if (main_genericstandalone_tx_init_tick) begin
				builder_a7_1000basex_gtptxinit_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_34 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_init_drpaddr = 5'd17;

// synthesis translate_off
reg dummy_d_35;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_init_drpdi <= 16'd0;
	if (main_genericstandalone_rx_init_drpmask) begin
		main_genericstandalone_rx_init_drpdi <= (main_genericstandalone_rx_init_drpvalue & 16'd63487);
	end else begin
		main_genericstandalone_rx_init_drpdi <= main_genericstandalone_rx_init_drpvalue;
	end
// synthesis translate_off
	dummy_d_35 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_36;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_init_drpen <= 1'd0;
	main_genericstandalone_rx_init_drpwe <= 1'd0;
	main_genericstandalone_rx_init_done <= 1'd0;
	main_genericstandalone_rx_init_rx_reset1 <= 1'd0;
	main_genericstandalone_rx_init_drpmask <= 1'd0;
	builder_a7_1000basex_gtprxinit_next_state <= 4'd0;
	main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value <= 16'd0;
	main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value_ce <= 1'd0;
	builder_a7_1000basex_gtprxinit_next_state <= builder_a7_1000basex_gtprxinit_state;
	case (builder_a7_1000basex_gtprxinit_state)
		1'd1: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			builder_a7_1000basex_gtprxinit_next_state <= 2'd2;
		end
		2'd2: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			main_genericstandalone_rx_init_drpen <= 1'd1;
			builder_a7_1000basex_gtprxinit_next_state <= 2'd3;
		end
		2'd3: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			if (main_genericstandalone_rx_init_drprdy) begin
				main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value <= main_genericstandalone_rx_init_drpdo;
				main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value_ce <= 1'd1;
				builder_a7_1000basex_gtprxinit_next_state <= 3'd4;
			end
		end
		3'd4: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			main_genericstandalone_rx_init_drpmask <= 1'd1;
			main_genericstandalone_rx_init_drpen <= 1'd1;
			main_genericstandalone_rx_init_drpwe <= 1'd1;
			builder_a7_1000basex_gtprxinit_next_state <= 3'd5;
		end
		3'd5: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			if (main_genericstandalone_rx_init_drprdy) begin
				builder_a7_1000basex_gtprxinit_next_state <= 3'd6;
			end
		end
		3'd6: begin
			if ((main_genericstandalone_rx_init_rx_pma_reset_done_r & (~main_genericstandalone_rx_init_rx_pma_reset_done1))) begin
				builder_a7_1000basex_gtprxinit_next_state <= 3'd7;
			end
		end
		3'd7: begin
			main_genericstandalone_rx_init_drpen <= 1'd1;
			main_genericstandalone_rx_init_drpwe <= 1'd1;
			builder_a7_1000basex_gtprxinit_next_state <= 4'd8;
		end
		4'd8: begin
			if (main_genericstandalone_rx_init_drprdy) begin
				builder_a7_1000basex_gtprxinit_next_state <= 4'd9;
			end
		end
		4'd9: begin
			main_genericstandalone_rx_init_done <= 1'd1;
			if (main_genericstandalone_rx_init_restart) begin
				builder_a7_1000basex_gtprxinit_next_state <= 1'd0;
			end
		end
		default: begin
			if (main_genericstandalone_rx_init_enable) begin
				builder_a7_1000basex_gtprxinit_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_36 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_o = (main_genericstandalone_toggle_o ^ main_genericstandalone_toggle_o_r);
assign main_genericstandalone_tx_cdc_sink_stb = main_genericstandalone_source_source_stb;
assign main_genericstandalone_source_source_ack = main_genericstandalone_tx_cdc_sink_ack;
assign main_genericstandalone_tx_cdc_sink_last = main_genericstandalone_source_source_last;
assign main_genericstandalone_tx_cdc_sink_eop = main_genericstandalone_source_source_eop;
assign main_genericstandalone_tx_cdc_sink_payload_data = main_genericstandalone_source_source_payload_data;
assign main_genericstandalone_tx_cdc_sink_payload_last_be = main_genericstandalone_source_source_payload_last_be;
assign main_genericstandalone_tx_cdc_sink_payload_error = main_genericstandalone_source_source_payload_error;
assign main_genericstandalone_sink_sink_stb = main_genericstandalone_rx_cdc_source_stb;
assign main_genericstandalone_rx_cdc_source_ack = main_genericstandalone_sink_sink_ack;
assign main_genericstandalone_sink_sink_last = main_genericstandalone_rx_cdc_source_last;
assign main_genericstandalone_sink_sink_eop = main_genericstandalone_rx_cdc_source_eop;
assign main_genericstandalone_sink_sink_payload_data = main_genericstandalone_rx_cdc_source_payload_data;
assign main_genericstandalone_sink_sink_payload_last_be = main_genericstandalone_rx_cdc_source_payload_last_be;
assign main_genericstandalone_sink_sink_payload_error = main_genericstandalone_rx_cdc_source_payload_error;
assign main_genericstandalone_ps_preamble_error_i = main_genericstandalone_preamble_checker_error;
assign main_genericstandalone_ps_crc_error_i = main_genericstandalone_crc32_checker_error;
assign main_genericstandalone_tx_converter_sink_sink_stb = main_genericstandalone_tx_cdc_source_stb;
assign main_genericstandalone_tx_cdc_source_ack = main_genericstandalone_tx_converter_sink_sink_ack;
assign main_genericstandalone_tx_converter_sink_sink_last = main_genericstandalone_tx_cdc_source_last;
assign main_genericstandalone_tx_converter_sink_sink_eop = main_genericstandalone_tx_cdc_source_eop;
assign main_genericstandalone_tx_converter_sink_sink_payload_data = main_genericstandalone_tx_cdc_source_payload_data;
assign main_genericstandalone_tx_converter_sink_sink_payload_last_be = main_genericstandalone_tx_cdc_source_payload_last_be;
assign main_genericstandalone_tx_converter_sink_sink_payload_error = main_genericstandalone_tx_cdc_source_payload_error;
assign main_genericstandalone_tx_last_be_sink_stb = main_genericstandalone_tx_converter_source_source_stb;
assign main_genericstandalone_tx_converter_source_source_ack = main_genericstandalone_tx_last_be_sink_ack;
assign main_genericstandalone_tx_last_be_sink_last = main_genericstandalone_tx_converter_source_source_last;
assign main_genericstandalone_tx_last_be_sink_eop = main_genericstandalone_tx_converter_source_source_eop;
assign main_genericstandalone_tx_last_be_sink_payload_data = main_genericstandalone_tx_converter_source_source_payload_data;
assign main_genericstandalone_tx_last_be_sink_payload_last_be = main_genericstandalone_tx_converter_source_source_payload_last_be;
assign main_genericstandalone_tx_last_be_sink_payload_error = main_genericstandalone_tx_converter_source_source_payload_error;
assign main_genericstandalone_padding_inserter_sink_stb = main_genericstandalone_tx_last_be_source_stb;
assign main_genericstandalone_tx_last_be_source_ack = main_genericstandalone_padding_inserter_sink_ack;
assign main_genericstandalone_padding_inserter_sink_last = main_genericstandalone_tx_last_be_source_last;
assign main_genericstandalone_padding_inserter_sink_eop = main_genericstandalone_tx_last_be_source_eop;
assign main_genericstandalone_padding_inserter_sink_payload_data = main_genericstandalone_tx_last_be_source_payload_data;
assign main_genericstandalone_padding_inserter_sink_payload_last_be = main_genericstandalone_tx_last_be_source_payload_last_be;
assign main_genericstandalone_padding_inserter_sink_payload_error = main_genericstandalone_tx_last_be_source_payload_error;
assign main_genericstandalone_crc32_inserter_sink_stb = main_genericstandalone_padding_inserter_source_stb;
assign main_genericstandalone_padding_inserter_source_ack = main_genericstandalone_crc32_inserter_sink_ack;
assign main_genericstandalone_crc32_inserter_sink_last = main_genericstandalone_padding_inserter_source_last;
assign main_genericstandalone_crc32_inserter_sink_eop = main_genericstandalone_padding_inserter_source_eop;
assign main_genericstandalone_crc32_inserter_sink_payload_data = main_genericstandalone_padding_inserter_source_payload_data;
assign main_genericstandalone_crc32_inserter_sink_payload_last_be = main_genericstandalone_padding_inserter_source_payload_last_be;
assign main_genericstandalone_crc32_inserter_sink_payload_error = main_genericstandalone_padding_inserter_source_payload_error;
assign main_genericstandalone_preamble_inserter_sink_stb = main_genericstandalone_crc32_inserter_source_stb;
assign main_genericstandalone_crc32_inserter_source_ack = main_genericstandalone_preamble_inserter_sink_ack;
assign main_genericstandalone_preamble_inserter_sink_last = main_genericstandalone_crc32_inserter_source_last;
assign main_genericstandalone_preamble_inserter_sink_eop = main_genericstandalone_crc32_inserter_source_eop;
assign main_genericstandalone_preamble_inserter_sink_payload_data = main_genericstandalone_crc32_inserter_source_payload_data;
assign main_genericstandalone_preamble_inserter_sink_payload_last_be = main_genericstandalone_crc32_inserter_source_payload_last_be;
assign main_genericstandalone_preamble_inserter_sink_payload_error = main_genericstandalone_crc32_inserter_source_payload_error;
assign main_genericstandalone_tx_gap_inserter_sink_stb = main_genericstandalone_preamble_inserter_source_stb;
assign main_genericstandalone_preamble_inserter_source_ack = main_genericstandalone_tx_gap_inserter_sink_ack;
assign main_genericstandalone_tx_gap_inserter_sink_last = main_genericstandalone_preamble_inserter_source_last;
assign main_genericstandalone_tx_gap_inserter_sink_eop = main_genericstandalone_preamble_inserter_source_eop;
assign main_genericstandalone_tx_gap_inserter_sink_payload_data = main_genericstandalone_preamble_inserter_source_payload_data;
assign main_genericstandalone_tx_gap_inserter_sink_payload_last_be = main_genericstandalone_preamble_inserter_source_payload_last_be;
assign main_genericstandalone_tx_gap_inserter_sink_payload_error = main_genericstandalone_preamble_inserter_source_payload_error;
assign main_genericstandalone_pcs_sink_stb = main_genericstandalone_tx_gap_inserter_source_stb;
assign main_genericstandalone_tx_gap_inserter_source_ack = main_genericstandalone_pcs_sink_ack;
assign main_genericstandalone_pcs_sink_last = main_genericstandalone_tx_gap_inserter_source_last;
assign main_genericstandalone_pcs_sink_eop = main_genericstandalone_tx_gap_inserter_source_eop;
assign main_genericstandalone_pcs_sink_payload_data = main_genericstandalone_tx_gap_inserter_source_payload_data;
assign main_genericstandalone_pcs_sink_payload_last_be = main_genericstandalone_tx_gap_inserter_source_payload_last_be;
assign main_genericstandalone_pcs_sink_payload_error = main_genericstandalone_tx_gap_inserter_source_payload_error;
assign main_genericstandalone_preamble_checker_sink_stb = main_genericstandalone_pcs_source_stb;
assign main_genericstandalone_pcs_source_ack = main_genericstandalone_preamble_checker_sink_ack;
assign main_genericstandalone_preamble_checker_sink_last = main_genericstandalone_pcs_source_last;
assign main_genericstandalone_preamble_checker_sink_eop = main_genericstandalone_pcs_source_eop;
assign main_genericstandalone_preamble_checker_sink_payload_data = main_genericstandalone_pcs_source_payload_data;
assign main_genericstandalone_preamble_checker_sink_payload_last_be = main_genericstandalone_pcs_source_payload_last_be;
assign main_genericstandalone_preamble_checker_sink_payload_error = main_genericstandalone_pcs_source_payload_error;
assign main_genericstandalone_crc32_checker_sink_sink_stb = main_genericstandalone_preamble_checker_source_stb;
assign main_genericstandalone_preamble_checker_source_ack = main_genericstandalone_crc32_checker_sink_sink_ack;
assign main_genericstandalone_crc32_checker_sink_sink_last = main_genericstandalone_preamble_checker_source_last;
assign main_genericstandalone_crc32_checker_sink_sink_eop = main_genericstandalone_preamble_checker_source_eop;
assign main_genericstandalone_crc32_checker_sink_sink_payload_data = main_genericstandalone_preamble_checker_source_payload_data;
assign main_genericstandalone_crc32_checker_sink_sink_payload_last_be = main_genericstandalone_preamble_checker_source_payload_last_be;
assign main_genericstandalone_crc32_checker_sink_sink_payload_error = main_genericstandalone_preamble_checker_source_payload_error;
assign main_genericstandalone_padding_checker_sink_stb = main_genericstandalone_crc32_checker_source_source_stb;
assign main_genericstandalone_crc32_checker_source_source_ack = main_genericstandalone_padding_checker_sink_ack;
assign main_genericstandalone_padding_checker_sink_last = main_genericstandalone_crc32_checker_source_source_last;
assign main_genericstandalone_padding_checker_sink_eop = main_genericstandalone_crc32_checker_source_source_eop;
assign main_genericstandalone_padding_checker_sink_payload_data = main_genericstandalone_crc32_checker_source_source_payload_data;
assign main_genericstandalone_padding_checker_sink_payload_last_be = main_genericstandalone_crc32_checker_source_source_payload_last_be;
assign main_genericstandalone_padding_checker_sink_payload_error = main_genericstandalone_crc32_checker_source_source_payload_error;
assign main_genericstandalone_rx_last_be_sink_stb = main_genericstandalone_padding_checker_source_stb;
assign main_genericstandalone_padding_checker_source_ack = main_genericstandalone_rx_last_be_sink_ack;
assign main_genericstandalone_rx_last_be_sink_last = main_genericstandalone_padding_checker_source_last;
assign main_genericstandalone_rx_last_be_sink_eop = main_genericstandalone_padding_checker_source_eop;
assign main_genericstandalone_rx_last_be_sink_payload_data = main_genericstandalone_padding_checker_source_payload_data;
assign main_genericstandalone_rx_last_be_sink_payload_last_be = main_genericstandalone_padding_checker_source_payload_last_be;
assign main_genericstandalone_rx_last_be_sink_payload_error = main_genericstandalone_padding_checker_source_payload_error;
assign main_genericstandalone_rx_converter_sink_sink_stb = main_genericstandalone_rx_last_be_source_stb;
assign main_genericstandalone_rx_last_be_source_ack = main_genericstandalone_rx_converter_sink_sink_ack;
assign main_genericstandalone_rx_converter_sink_sink_last = main_genericstandalone_rx_last_be_source_last;
assign main_genericstandalone_rx_converter_sink_sink_eop = main_genericstandalone_rx_last_be_source_eop;
assign main_genericstandalone_rx_converter_sink_sink_payload_data = main_genericstandalone_rx_last_be_source_payload_data;
assign main_genericstandalone_rx_converter_sink_sink_payload_last_be = main_genericstandalone_rx_last_be_source_payload_last_be;
assign main_genericstandalone_rx_converter_sink_sink_payload_error = main_genericstandalone_rx_last_be_source_payload_error;
assign main_genericstandalone_rx_cdc_sink_stb = main_genericstandalone_rx_converter_source_source_stb;
assign main_genericstandalone_rx_converter_source_source_ack = main_genericstandalone_rx_cdc_sink_ack;
assign main_genericstandalone_rx_cdc_sink_last = main_genericstandalone_rx_converter_source_source_last;
assign main_genericstandalone_rx_cdc_sink_eop = main_genericstandalone_rx_converter_source_source_eop;
assign main_genericstandalone_rx_cdc_sink_payload_data = main_genericstandalone_rx_converter_source_source_payload_data;
assign main_genericstandalone_rx_cdc_sink_payload_last_be = main_genericstandalone_rx_converter_source_source_payload_last_be;
assign main_genericstandalone_rx_cdc_sink_payload_error = main_genericstandalone_rx_converter_source_source_payload_error;

// synthesis translate_off
reg dummy_d_37;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_gap_inserter_sink_ack <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_stb <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_last <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_eop <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_payload_data <= 8'd0;
	main_genericstandalone_tx_gap_inserter_source_payload_last_be <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_payload_error <= 1'd0;
	main_genericstandalone_tx_gap_inserter_counter_reset <= 1'd0;
	main_genericstandalone_tx_gap_inserter_counter_ce <= 1'd0;
	builder_liteethmacgap_next_state <= 1'd0;
	builder_liteethmacgap_next_state <= builder_liteethmacgap_state;
	case (builder_liteethmacgap_state)
		1'd1: begin
			main_genericstandalone_tx_gap_inserter_counter_ce <= 1'd1;
			if ((main_genericstandalone_tx_gap_inserter_counter == 4'd11)) begin
				builder_liteethmacgap_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_tx_gap_inserter_counter_reset <= 1'd1;
			main_genericstandalone_tx_gap_inserter_source_stb <= main_genericstandalone_tx_gap_inserter_sink_stb;
			main_genericstandalone_tx_gap_inserter_sink_ack <= main_genericstandalone_tx_gap_inserter_source_ack;
			main_genericstandalone_tx_gap_inserter_source_last <= main_genericstandalone_tx_gap_inserter_sink_last;
			main_genericstandalone_tx_gap_inserter_source_eop <= main_genericstandalone_tx_gap_inserter_sink_eop;
			main_genericstandalone_tx_gap_inserter_source_payload_data <= main_genericstandalone_tx_gap_inserter_sink_payload_data;
			main_genericstandalone_tx_gap_inserter_source_payload_last_be <= main_genericstandalone_tx_gap_inserter_sink_payload_last_be;
			main_genericstandalone_tx_gap_inserter_source_payload_error <= main_genericstandalone_tx_gap_inserter_sink_payload_error;
			if (((main_genericstandalone_tx_gap_inserter_sink_stb & main_genericstandalone_tx_gap_inserter_sink_eop) & main_genericstandalone_tx_gap_inserter_sink_ack)) begin
				builder_liteethmacgap_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_37 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_preamble_inserter_source_payload_last_be = main_genericstandalone_preamble_inserter_sink_payload_last_be;

// synthesis translate_off
reg dummy_d_38;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_preamble_inserter_sink_ack <= 1'd0;
	main_genericstandalone_preamble_inserter_source_stb <= 1'd0;
	main_genericstandalone_preamble_inserter_source_last <= 1'd0;
	main_genericstandalone_preamble_inserter_source_eop <= 1'd0;
	main_genericstandalone_preamble_inserter_source_payload_data <= 8'd0;
	main_genericstandalone_preamble_inserter_source_payload_error <= 1'd0;
	main_genericstandalone_preamble_inserter_clr_cnt <= 1'd0;
	main_genericstandalone_preamble_inserter_inc_cnt <= 1'd0;
	builder_liteethmacpreambleinserter_next_state <= 2'd0;
	main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_sink_payload_data;
	builder_liteethmacpreambleinserter_next_state <= builder_liteethmacpreambleinserter_state;
	case (builder_liteethmacpreambleinserter_state)
		1'd1: begin
			main_genericstandalone_preamble_inserter_source_stb <= 1'd1;
			case (main_genericstandalone_preamble_inserter_cnt)
				1'd0: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[7:0];
				end
				1'd1: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[15:8];
				end
				2'd2: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[23:16];
				end
				2'd3: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[31:24];
				end
				3'd4: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[39:32];
				end
				3'd5: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[47:40];
				end
				3'd6: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[55:48];
				end
				default: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[63:56];
				end
			endcase
			if ((main_genericstandalone_preamble_inserter_cnt == 3'd7)) begin
				if (main_genericstandalone_preamble_inserter_source_ack) begin
					builder_liteethmacpreambleinserter_next_state <= 2'd2;
				end
			end else begin
				main_genericstandalone_preamble_inserter_inc_cnt <= main_genericstandalone_preamble_inserter_source_ack;
			end
		end
		2'd2: begin
			main_genericstandalone_preamble_inserter_source_stb <= main_genericstandalone_preamble_inserter_sink_stb;
			main_genericstandalone_preamble_inserter_sink_ack <= main_genericstandalone_preamble_inserter_source_ack;
			main_genericstandalone_preamble_inserter_source_last <= main_genericstandalone_preamble_inserter_sink_last;
			main_genericstandalone_preamble_inserter_source_eop <= main_genericstandalone_preamble_inserter_sink_eop;
			main_genericstandalone_preamble_inserter_source_payload_error <= main_genericstandalone_preamble_inserter_sink_payload_error;
			if (((main_genericstandalone_preamble_inserter_sink_stb & main_genericstandalone_preamble_inserter_sink_eop) & main_genericstandalone_preamble_inserter_source_ack)) begin
				builder_liteethmacpreambleinserter_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_preamble_inserter_sink_ack <= 1'd1;
			main_genericstandalone_preamble_inserter_clr_cnt <= 1'd1;
			if (main_genericstandalone_preamble_inserter_sink_stb) begin
				main_genericstandalone_preamble_inserter_sink_ack <= 1'd0;
				builder_liteethmacpreambleinserter_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_38 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_preamble_checker_source_payload_data = main_genericstandalone_preamble_checker_sink_payload_data;
assign main_genericstandalone_preamble_checker_source_payload_last_be = main_genericstandalone_preamble_checker_sink_payload_last_be;

// synthesis translate_off
reg dummy_d_39;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_preamble_checker_sink_ack <= 1'd0;
	main_genericstandalone_preamble_checker_source_stb <= 1'd0;
	main_genericstandalone_preamble_checker_source_last <= 1'd0;
	main_genericstandalone_preamble_checker_source_eop <= 1'd0;
	main_genericstandalone_preamble_checker_source_payload_error <= 1'd0;
	main_genericstandalone_preamble_checker_error <= 1'd0;
	builder_liteethmacpreamblechecker_next_state <= 1'd0;
	builder_liteethmacpreamblechecker_next_state <= builder_liteethmacpreamblechecker_state;
	case (builder_liteethmacpreamblechecker_state)
		1'd1: begin
			main_genericstandalone_preamble_checker_source_stb <= main_genericstandalone_preamble_checker_sink_stb;
			main_genericstandalone_preamble_checker_sink_ack <= main_genericstandalone_preamble_checker_source_ack;
			main_genericstandalone_preamble_checker_source_last <= main_genericstandalone_preamble_checker_sink_last;
			main_genericstandalone_preamble_checker_source_eop <= main_genericstandalone_preamble_checker_sink_eop;
			main_genericstandalone_preamble_checker_source_payload_error <= main_genericstandalone_preamble_checker_sink_payload_error;
			if (((main_genericstandalone_preamble_checker_source_stb & main_genericstandalone_preamble_checker_source_eop) & main_genericstandalone_preamble_checker_source_ack)) begin
				builder_liteethmacpreamblechecker_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_preamble_checker_sink_ack <= 1'd1;
			if (((main_genericstandalone_preamble_checker_sink_stb & (~main_genericstandalone_preamble_checker_sink_eop)) & (main_genericstandalone_preamble_checker_sink_payload_data == 8'd213))) begin
				builder_liteethmacpreamblechecker_next_state <= 1'd1;
			end
			if ((main_genericstandalone_preamble_checker_sink_stb & main_genericstandalone_preamble_checker_sink_eop)) begin
				main_genericstandalone_preamble_checker_error <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_39 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_inserter_cnt_done = (main_genericstandalone_crc32_inserter_cnt == 1'd0);
assign main_genericstandalone_crc32_inserter_data1 = main_genericstandalone_crc32_inserter_data0;
assign main_genericstandalone_crc32_inserter_last = main_genericstandalone_crc32_inserter_reg;
assign main_genericstandalone_crc32_inserter_value = (~{main_genericstandalone_crc32_inserter_reg[0], main_genericstandalone_crc32_inserter_reg[1], main_genericstandalone_crc32_inserter_reg[2], main_genericstandalone_crc32_inserter_reg[3], main_genericstandalone_crc32_inserter_reg[4], main_genericstandalone_crc32_inserter_reg[5], main_genericstandalone_crc32_inserter_reg[6], main_genericstandalone_crc32_inserter_reg[7], main_genericstandalone_crc32_inserter_reg[8], main_genericstandalone_crc32_inserter_reg[9], main_genericstandalone_crc32_inserter_reg[10], main_genericstandalone_crc32_inserter_reg[11], main_genericstandalone_crc32_inserter_reg[12], main_genericstandalone_crc32_inserter_reg[13], main_genericstandalone_crc32_inserter_reg[14], main_genericstandalone_crc32_inserter_reg[15], main_genericstandalone_crc32_inserter_reg[16], main_genericstandalone_crc32_inserter_reg[17], main_genericstandalone_crc32_inserter_reg[18], main_genericstandalone_crc32_inserter_reg[19], main_genericstandalone_crc32_inserter_reg[20], main_genericstandalone_crc32_inserter_reg[21], main_genericstandalone_crc32_inserter_reg[22], main_genericstandalone_crc32_inserter_reg[23], main_genericstandalone_crc32_inserter_reg[24], main_genericstandalone_crc32_inserter_reg[25], main_genericstandalone_crc32_inserter_reg[26], main_genericstandalone_crc32_inserter_reg[27], main_genericstandalone_crc32_inserter_reg[28], main_genericstandalone_crc32_inserter_reg[29], main_genericstandalone_crc32_inserter_reg[30], main_genericstandalone_crc32_inserter_reg[31]});
assign main_genericstandalone_crc32_inserter_error = (main_genericstandalone_crc32_inserter_next != 32'd3338984827);

// synthesis translate_off
reg dummy_d_40;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_inserter_next <= 32'd0;
	main_genericstandalone_crc32_inserter_next[0] <= (((main_genericstandalone_crc32_inserter_last[24] ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[1] <= (((((((main_genericstandalone_crc32_inserter_last[25] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[2] <= (((((((((main_genericstandalone_crc32_inserter_last[26] ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[3] <= (((((((main_genericstandalone_crc32_inserter_last[27] ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[4] <= (((((((((main_genericstandalone_crc32_inserter_last[28] ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[5] <= (((((((((((((main_genericstandalone_crc32_inserter_last[29] ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[6] <= (((((((((((main_genericstandalone_crc32_inserter_last[30] ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[7] <= (((((((((main_genericstandalone_crc32_inserter_last[31] ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[8] <= ((((((((main_genericstandalone_crc32_inserter_last[0] ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[9] <= ((((((((main_genericstandalone_crc32_inserter_last[1] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[10] <= ((((((((main_genericstandalone_crc32_inserter_last[2] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[11] <= ((((((((main_genericstandalone_crc32_inserter_last[3] ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[12] <= ((((((((((((main_genericstandalone_crc32_inserter_last[4] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[13] <= ((((((((((((main_genericstandalone_crc32_inserter_last[5] ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[14] <= ((((((((((main_genericstandalone_crc32_inserter_last[6] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]);
	main_genericstandalone_crc32_inserter_next[15] <= ((((((((main_genericstandalone_crc32_inserter_last[7] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]);
	main_genericstandalone_crc32_inserter_next[16] <= ((((((main_genericstandalone_crc32_inserter_last[8] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[17] <= ((((((main_genericstandalone_crc32_inserter_last[9] ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[18] <= ((((((main_genericstandalone_crc32_inserter_last[10] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]);
	main_genericstandalone_crc32_inserter_next[19] <= ((((main_genericstandalone_crc32_inserter_last[11] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]);
	main_genericstandalone_crc32_inserter_next[20] <= ((main_genericstandalone_crc32_inserter_last[12] ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]);
	main_genericstandalone_crc32_inserter_next[21] <= ((main_genericstandalone_crc32_inserter_last[13] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]);
	main_genericstandalone_crc32_inserter_next[22] <= ((main_genericstandalone_crc32_inserter_last[14] ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[23] <= ((((((main_genericstandalone_crc32_inserter_last[15] ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[24] <= ((((((main_genericstandalone_crc32_inserter_last[16] ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[25] <= ((((main_genericstandalone_crc32_inserter_last[17] ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]);
	main_genericstandalone_crc32_inserter_next[26] <= ((((((((main_genericstandalone_crc32_inserter_last[18] ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[27] <= ((((((((main_genericstandalone_crc32_inserter_last[19] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[28] <= ((((((main_genericstandalone_crc32_inserter_last[20] ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]);
	main_genericstandalone_crc32_inserter_next[29] <= ((((((main_genericstandalone_crc32_inserter_last[21] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]);
	main_genericstandalone_crc32_inserter_next[30] <= ((((main_genericstandalone_crc32_inserter_last[22] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]);
	main_genericstandalone_crc32_inserter_next[31] <= ((main_genericstandalone_crc32_inserter_last[23] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]);
// synthesis translate_off
	dummy_d_40 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_41;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_inserter_sink_ack <= 1'd0;
	main_genericstandalone_crc32_inserter_source_stb <= 1'd0;
	main_genericstandalone_crc32_inserter_source_last <= 1'd0;
	main_genericstandalone_crc32_inserter_source_eop <= 1'd0;
	main_genericstandalone_crc32_inserter_source_payload_data <= 8'd0;
	main_genericstandalone_crc32_inserter_source_payload_last_be <= 1'd0;
	main_genericstandalone_crc32_inserter_source_payload_error <= 1'd0;
	main_genericstandalone_crc32_inserter_data0 <= 8'd0;
	main_genericstandalone_crc32_inserter_ce <= 1'd0;
	main_genericstandalone_crc32_inserter_reset <= 1'd0;
	main_genericstandalone_crc32_inserter_is_ongoing0 <= 1'd0;
	main_genericstandalone_crc32_inserter_is_ongoing1 <= 1'd0;
	builder_liteethmaccrc32inserter_next_state <= 2'd0;
	builder_liteethmaccrc32inserter_next_state <= builder_liteethmaccrc32inserter_state;
	case (builder_liteethmaccrc32inserter_state)
		1'd1: begin
			main_genericstandalone_crc32_inserter_ce <= (main_genericstandalone_crc32_inserter_sink_stb & main_genericstandalone_crc32_inserter_source_ack);
			main_genericstandalone_crc32_inserter_data0 <= main_genericstandalone_crc32_inserter_sink_payload_data;
			main_genericstandalone_crc32_inserter_source_stb <= main_genericstandalone_crc32_inserter_sink_stb;
			main_genericstandalone_crc32_inserter_sink_ack <= main_genericstandalone_crc32_inserter_source_ack;
			main_genericstandalone_crc32_inserter_source_last <= main_genericstandalone_crc32_inserter_sink_last;
			main_genericstandalone_crc32_inserter_source_eop <= main_genericstandalone_crc32_inserter_sink_eop;
			main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_sink_payload_data;
			main_genericstandalone_crc32_inserter_source_payload_last_be <= main_genericstandalone_crc32_inserter_sink_payload_last_be;
			main_genericstandalone_crc32_inserter_source_payload_error <= main_genericstandalone_crc32_inserter_sink_payload_error;
			main_genericstandalone_crc32_inserter_source_eop <= 1'd0;
			if (((main_genericstandalone_crc32_inserter_sink_stb & main_genericstandalone_crc32_inserter_sink_eop) & main_genericstandalone_crc32_inserter_source_ack)) begin
				builder_liteethmaccrc32inserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_genericstandalone_crc32_inserter_source_stb <= 1'd1;
			case (main_genericstandalone_crc32_inserter_cnt)
				1'd0: begin
					main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_value[31:24];
				end
				1'd1: begin
					main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_value[23:16];
				end
				2'd2: begin
					main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_value[15:8];
				end
				default: begin
					main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_value[7:0];
				end
			endcase
			if (main_genericstandalone_crc32_inserter_cnt_done) begin
				main_genericstandalone_crc32_inserter_source_eop <= 1'd1;
				if (main_genericstandalone_crc32_inserter_source_ack) begin
					builder_liteethmaccrc32inserter_next_state <= 1'd0;
				end
			end
			main_genericstandalone_crc32_inserter_is_ongoing1 <= 1'd1;
		end
		default: begin
			main_genericstandalone_crc32_inserter_reset <= 1'd1;
			main_genericstandalone_crc32_inserter_sink_ack <= 1'd1;
			if (main_genericstandalone_crc32_inserter_sink_stb) begin
				main_genericstandalone_crc32_inserter_sink_ack <= 1'd0;
				builder_liteethmaccrc32inserter_next_state <= 1'd1;
			end
			main_genericstandalone_crc32_inserter_is_ongoing0 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_41 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_fifo_full = (main_genericstandalone_crc32_checker_syncfifo_level == 3'd4);
assign main_genericstandalone_crc32_checker_fifo_in = (main_genericstandalone_crc32_checker_sink_sink_stb & ((~main_genericstandalone_crc32_checker_fifo_full) | main_genericstandalone_crc32_checker_fifo_out));
assign main_genericstandalone_crc32_checker_fifo_out = (main_genericstandalone_crc32_checker_source_source_stb & main_genericstandalone_crc32_checker_source_source_ack);
assign main_genericstandalone_crc32_checker_syncfifo_sink_last = main_genericstandalone_crc32_checker_sink_sink_last;
assign main_genericstandalone_crc32_checker_syncfifo_sink_eop = main_genericstandalone_crc32_checker_sink_sink_eop;
assign main_genericstandalone_crc32_checker_syncfifo_sink_payload_data = main_genericstandalone_crc32_checker_sink_sink_payload_data;
assign main_genericstandalone_crc32_checker_syncfifo_sink_payload_last_be = main_genericstandalone_crc32_checker_sink_sink_payload_last_be;
assign main_genericstandalone_crc32_checker_syncfifo_sink_payload_error = main_genericstandalone_crc32_checker_sink_sink_payload_error;

// synthesis translate_off
reg dummy_d_42;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_syncfifo_sink_stb <= 1'd0;
	main_genericstandalone_crc32_checker_syncfifo_sink_stb <= main_genericstandalone_crc32_checker_sink_sink_stb;
	main_genericstandalone_crc32_checker_syncfifo_sink_stb <= main_genericstandalone_crc32_checker_fifo_in;
// synthesis translate_off
	dummy_d_42 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_43;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_sink_sink_ack <= 1'd0;
	main_genericstandalone_crc32_checker_sink_sink_ack <= main_genericstandalone_crc32_checker_syncfifo_sink_ack;
	main_genericstandalone_crc32_checker_sink_sink_ack <= main_genericstandalone_crc32_checker_fifo_in;
// synthesis translate_off
	dummy_d_43 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_source_source_stb = (main_genericstandalone_crc32_checker_sink_sink_stb & main_genericstandalone_crc32_checker_fifo_full);
assign main_genericstandalone_crc32_checker_source_source_eop = main_genericstandalone_crc32_checker_sink_sink_eop;
assign main_genericstandalone_crc32_checker_syncfifo_source_ack = main_genericstandalone_crc32_checker_fifo_out;
assign main_genericstandalone_crc32_checker_source_source_payload_data = main_genericstandalone_crc32_checker_syncfifo_source_payload_data;
assign main_genericstandalone_crc32_checker_source_source_payload_last_be = main_genericstandalone_crc32_checker_syncfifo_source_payload_last_be;

// synthesis translate_off
reg dummy_d_44;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_source_source_payload_error <= 1'd0;
	main_genericstandalone_crc32_checker_source_source_payload_error <= main_genericstandalone_crc32_checker_syncfifo_source_payload_error;
	main_genericstandalone_crc32_checker_source_source_payload_error <= (main_genericstandalone_crc32_checker_sink_sink_payload_error | main_genericstandalone_crc32_checker_crc_error);
// synthesis translate_off
	dummy_d_44 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_error = ((main_genericstandalone_crc32_checker_source_source_stb & main_genericstandalone_crc32_checker_source_source_eop) & main_genericstandalone_crc32_checker_crc_error);
assign main_genericstandalone_crc32_checker_crc_data0 = main_genericstandalone_crc32_checker_sink_sink_payload_data;
assign main_genericstandalone_crc32_checker_crc_data1 = main_genericstandalone_crc32_checker_crc_data0;
assign main_genericstandalone_crc32_checker_crc_last = main_genericstandalone_crc32_checker_crc_reg;
assign main_genericstandalone_crc32_checker_crc_value = (~{main_genericstandalone_crc32_checker_crc_reg[0], main_genericstandalone_crc32_checker_crc_reg[1], main_genericstandalone_crc32_checker_crc_reg[2], main_genericstandalone_crc32_checker_crc_reg[3], main_genericstandalone_crc32_checker_crc_reg[4], main_genericstandalone_crc32_checker_crc_reg[5], main_genericstandalone_crc32_checker_crc_reg[6], main_genericstandalone_crc32_checker_crc_reg[7], main_genericstandalone_crc32_checker_crc_reg[8], main_genericstandalone_crc32_checker_crc_reg[9], main_genericstandalone_crc32_checker_crc_reg[10], main_genericstandalone_crc32_checker_crc_reg[11], main_genericstandalone_crc32_checker_crc_reg[12], main_genericstandalone_crc32_checker_crc_reg[13], main_genericstandalone_crc32_checker_crc_reg[14], main_genericstandalone_crc32_checker_crc_reg[15], main_genericstandalone_crc32_checker_crc_reg[16], main_genericstandalone_crc32_checker_crc_reg[17], main_genericstandalone_crc32_checker_crc_reg[18], main_genericstandalone_crc32_checker_crc_reg[19], main_genericstandalone_crc32_checker_crc_reg[20], main_genericstandalone_crc32_checker_crc_reg[21], main_genericstandalone_crc32_checker_crc_reg[22], main_genericstandalone_crc32_checker_crc_reg[23], main_genericstandalone_crc32_checker_crc_reg[24], main_genericstandalone_crc32_checker_crc_reg[25], main_genericstandalone_crc32_checker_crc_reg[26], main_genericstandalone_crc32_checker_crc_reg[27], main_genericstandalone_crc32_checker_crc_reg[28], main_genericstandalone_crc32_checker_crc_reg[29], main_genericstandalone_crc32_checker_crc_reg[30], main_genericstandalone_crc32_checker_crc_reg[31]});
assign main_genericstandalone_crc32_checker_crc_error = (main_genericstandalone_crc32_checker_crc_next != 32'd3338984827);

// synthesis translate_off
reg dummy_d_45;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_crc_next <= 32'd0;
	main_genericstandalone_crc32_checker_crc_next[0] <= (((main_genericstandalone_crc32_checker_crc_last[24] ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[1] <= (((((((main_genericstandalone_crc32_checker_crc_last[25] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[2] <= (((((((((main_genericstandalone_crc32_checker_crc_last[26] ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[3] <= (((((((main_genericstandalone_crc32_checker_crc_last[27] ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[4] <= (((((((((main_genericstandalone_crc32_checker_crc_last[28] ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[5] <= (((((((((((((main_genericstandalone_crc32_checker_crc_last[29] ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[6] <= (((((((((((main_genericstandalone_crc32_checker_crc_last[30] ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[7] <= (((((((((main_genericstandalone_crc32_checker_crc_last[31] ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[8] <= ((((((((main_genericstandalone_crc32_checker_crc_last[0] ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[9] <= ((((((((main_genericstandalone_crc32_checker_crc_last[1] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[10] <= ((((((((main_genericstandalone_crc32_checker_crc_last[2] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[11] <= ((((((((main_genericstandalone_crc32_checker_crc_last[3] ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[12] <= ((((((((((((main_genericstandalone_crc32_checker_crc_last[4] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[13] <= ((((((((((((main_genericstandalone_crc32_checker_crc_last[5] ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[14] <= ((((((((((main_genericstandalone_crc32_checker_crc_last[6] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]);
	main_genericstandalone_crc32_checker_crc_next[15] <= ((((((((main_genericstandalone_crc32_checker_crc_last[7] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]);
	main_genericstandalone_crc32_checker_crc_next[16] <= ((((((main_genericstandalone_crc32_checker_crc_last[8] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[17] <= ((((((main_genericstandalone_crc32_checker_crc_last[9] ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[18] <= ((((((main_genericstandalone_crc32_checker_crc_last[10] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]);
	main_genericstandalone_crc32_checker_crc_next[19] <= ((((main_genericstandalone_crc32_checker_crc_last[11] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]);
	main_genericstandalone_crc32_checker_crc_next[20] <= ((main_genericstandalone_crc32_checker_crc_last[12] ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]);
	main_genericstandalone_crc32_checker_crc_next[21] <= ((main_genericstandalone_crc32_checker_crc_last[13] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]);
	main_genericstandalone_crc32_checker_crc_next[22] <= ((main_genericstandalone_crc32_checker_crc_last[14] ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[23] <= ((((((main_genericstandalone_crc32_checker_crc_last[15] ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[24] <= ((((((main_genericstandalone_crc32_checker_crc_last[16] ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[25] <= ((((main_genericstandalone_crc32_checker_crc_last[17] ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]);
	main_genericstandalone_crc32_checker_crc_next[26] <= ((((((((main_genericstandalone_crc32_checker_crc_last[18] ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[27] <= ((((((((main_genericstandalone_crc32_checker_crc_last[19] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[28] <= ((((((main_genericstandalone_crc32_checker_crc_last[20] ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]);
	main_genericstandalone_crc32_checker_crc_next[29] <= ((((((main_genericstandalone_crc32_checker_crc_last[21] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]);
	main_genericstandalone_crc32_checker_crc_next[30] <= ((((main_genericstandalone_crc32_checker_crc_last[22] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]);
	main_genericstandalone_crc32_checker_crc_next[31] <= ((main_genericstandalone_crc32_checker_crc_last[23] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]);
// synthesis translate_off
	dummy_d_45 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_din = {main_genericstandalone_crc32_checker_syncfifo_fifo_in_eop, main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_error, main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_last_be, main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_data};
assign {main_genericstandalone_crc32_checker_syncfifo_fifo_out_eop, main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_error, main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_last_be, main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_data} = main_genericstandalone_crc32_checker_syncfifo_syncfifo_dout;
assign main_genericstandalone_crc32_checker_syncfifo_sink_ack = main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable;
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_we = main_genericstandalone_crc32_checker_syncfifo_sink_stb;
assign main_genericstandalone_crc32_checker_syncfifo_fifo_in_eop = main_genericstandalone_crc32_checker_syncfifo_sink_eop;
assign main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_data = main_genericstandalone_crc32_checker_syncfifo_sink_payload_data;
assign main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_last_be = main_genericstandalone_crc32_checker_syncfifo_sink_payload_last_be;
assign main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_error = main_genericstandalone_crc32_checker_syncfifo_sink_payload_error;
assign main_genericstandalone_crc32_checker_syncfifo_source_stb = main_genericstandalone_crc32_checker_syncfifo_syncfifo_readable;
assign main_genericstandalone_crc32_checker_syncfifo_source_eop = main_genericstandalone_crc32_checker_syncfifo_fifo_out_eop;
assign main_genericstandalone_crc32_checker_syncfifo_source_payload_data = main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_data;
assign main_genericstandalone_crc32_checker_syncfifo_source_payload_last_be = main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_last_be;
assign main_genericstandalone_crc32_checker_syncfifo_source_payload_error = main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_error;
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_re = main_genericstandalone_crc32_checker_syncfifo_source_ack;

// synthesis translate_off
reg dummy_d_46;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_syncfifo_wrport_adr <= 3'd0;
	if (main_genericstandalone_crc32_checker_syncfifo_replace) begin
		main_genericstandalone_crc32_checker_syncfifo_wrport_adr <= (main_genericstandalone_crc32_checker_syncfifo_produce - 1'd1);
	end else begin
		main_genericstandalone_crc32_checker_syncfifo_wrport_adr <= main_genericstandalone_crc32_checker_syncfifo_produce;
	end
// synthesis translate_off
	dummy_d_46 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_syncfifo_wrport_dat_w = main_genericstandalone_crc32_checker_syncfifo_syncfifo_din;
assign main_genericstandalone_crc32_checker_syncfifo_wrport_we = (main_genericstandalone_crc32_checker_syncfifo_syncfifo_we & (main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable | main_genericstandalone_crc32_checker_syncfifo_replace));
assign main_genericstandalone_crc32_checker_syncfifo_do_read = (main_genericstandalone_crc32_checker_syncfifo_syncfifo_readable & main_genericstandalone_crc32_checker_syncfifo_syncfifo_re);
assign main_genericstandalone_crc32_checker_syncfifo_rdport_adr = main_genericstandalone_crc32_checker_syncfifo_consume;
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_dout = main_genericstandalone_crc32_checker_syncfifo_rdport_dat_r;
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable = (main_genericstandalone_crc32_checker_syncfifo_level != 3'd5);
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_readable = (main_genericstandalone_crc32_checker_syncfifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_47;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_crc_ce <= 1'd0;
	main_genericstandalone_crc32_checker_crc_reset <= 1'd0;
	main_genericstandalone_crc32_checker_fifo_reset <= 1'd0;
	builder_liteethmaccrc32checker_next_state <= 2'd0;
	builder_liteethmaccrc32checker_next_state <= builder_liteethmaccrc32checker_state;
	case (builder_liteethmaccrc32checker_state)
		1'd1: begin
			if ((main_genericstandalone_crc32_checker_sink_sink_stb & main_genericstandalone_crc32_checker_sink_sink_ack)) begin
				main_genericstandalone_crc32_checker_crc_ce <= 1'd1;
				builder_liteethmaccrc32checker_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((main_genericstandalone_crc32_checker_sink_sink_stb & main_genericstandalone_crc32_checker_sink_sink_ack)) begin
				main_genericstandalone_crc32_checker_crc_ce <= 1'd1;
				if (main_genericstandalone_crc32_checker_sink_sink_eop) begin
					builder_liteethmaccrc32checker_next_state <= 1'd0;
				end
			end
		end
		default: begin
			main_genericstandalone_crc32_checker_crc_reset <= 1'd1;
			main_genericstandalone_crc32_checker_fifo_reset <= 1'd1;
			builder_liteethmaccrc32checker_next_state <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_47 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_ps_preamble_error_o = (main_genericstandalone_ps_preamble_error_toggle_o ^ main_genericstandalone_ps_preamble_error_toggle_o_r);
assign main_genericstandalone_ps_crc_error_o = (main_genericstandalone_ps_crc_error_toggle_o ^ main_genericstandalone_ps_crc_error_toggle_o_r);
assign main_genericstandalone_padding_inserter_counter_done = (main_genericstandalone_padding_inserter_counter >= 6'd59);

// synthesis translate_off
reg dummy_d_48;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_padding_inserter_sink_ack <= 1'd0;
	main_genericstandalone_padding_inserter_source_stb <= 1'd0;
	main_genericstandalone_padding_inserter_source_last <= 1'd0;
	main_genericstandalone_padding_inserter_source_eop <= 1'd0;
	main_genericstandalone_padding_inserter_source_payload_data <= 8'd0;
	main_genericstandalone_padding_inserter_source_payload_last_be <= 1'd0;
	main_genericstandalone_padding_inserter_source_payload_error <= 1'd0;
	main_genericstandalone_padding_inserter_counter_reset <= 1'd0;
	main_genericstandalone_padding_inserter_counter_ce <= 1'd0;
	builder_liteethmacpaddinginserter_next_state <= 1'd0;
	builder_liteethmacpaddinginserter_next_state <= builder_liteethmacpaddinginserter_state;
	case (builder_liteethmacpaddinginserter_state)
		1'd1: begin
			main_genericstandalone_padding_inserter_source_stb <= 1'd1;
			main_genericstandalone_padding_inserter_source_eop <= main_genericstandalone_padding_inserter_counter_done;
			main_genericstandalone_padding_inserter_source_payload_data <= 1'd0;
			if ((main_genericstandalone_padding_inserter_source_stb & main_genericstandalone_padding_inserter_source_ack)) begin
				main_genericstandalone_padding_inserter_counter_ce <= 1'd1;
				if (main_genericstandalone_padding_inserter_counter_done) begin
					main_genericstandalone_padding_inserter_counter_reset <= 1'd1;
					builder_liteethmacpaddinginserter_next_state <= 1'd0;
				end
			end
		end
		default: begin
			main_genericstandalone_padding_inserter_source_stb <= main_genericstandalone_padding_inserter_sink_stb;
			main_genericstandalone_padding_inserter_sink_ack <= main_genericstandalone_padding_inserter_source_ack;
			main_genericstandalone_padding_inserter_source_last <= main_genericstandalone_padding_inserter_sink_last;
			main_genericstandalone_padding_inserter_source_eop <= main_genericstandalone_padding_inserter_sink_eop;
			main_genericstandalone_padding_inserter_source_payload_data <= main_genericstandalone_padding_inserter_sink_payload_data;
			main_genericstandalone_padding_inserter_source_payload_last_be <= main_genericstandalone_padding_inserter_sink_payload_last_be;
			main_genericstandalone_padding_inserter_source_payload_error <= main_genericstandalone_padding_inserter_sink_payload_error;
			if ((main_genericstandalone_padding_inserter_source_stb & main_genericstandalone_padding_inserter_source_ack)) begin
				main_genericstandalone_padding_inserter_counter_ce <= 1'd1;
				if (main_genericstandalone_padding_inserter_sink_eop) begin
					if ((~main_genericstandalone_padding_inserter_counter_done)) begin
						main_genericstandalone_padding_inserter_source_eop <= 1'd0;
						builder_liteethmacpaddinginserter_next_state <= 1'd1;
					end else begin
						main_genericstandalone_padding_inserter_counter_reset <= 1'd1;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_48 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_padding_checker_source_stb = main_genericstandalone_padding_checker_sink_stb;
assign main_genericstandalone_padding_checker_sink_ack = main_genericstandalone_padding_checker_source_ack;
assign main_genericstandalone_padding_checker_source_last = main_genericstandalone_padding_checker_sink_last;
assign main_genericstandalone_padding_checker_source_eop = main_genericstandalone_padding_checker_sink_eop;
assign main_genericstandalone_padding_checker_source_payload_data = main_genericstandalone_padding_checker_sink_payload_data;
assign main_genericstandalone_padding_checker_source_payload_last_be = main_genericstandalone_padding_checker_sink_payload_last_be;
assign main_genericstandalone_padding_checker_source_payload_error = main_genericstandalone_padding_checker_sink_payload_error;
assign main_genericstandalone_tx_last_be_source_stb = (main_genericstandalone_tx_last_be_sink_stb & main_genericstandalone_tx_last_be_ongoing);
assign main_genericstandalone_tx_last_be_source_eop = main_genericstandalone_tx_last_be_sink_payload_last_be;
assign main_genericstandalone_tx_last_be_source_payload_data = main_genericstandalone_tx_last_be_sink_payload_data;
assign main_genericstandalone_tx_last_be_sink_ack = main_genericstandalone_tx_last_be_source_ack;
assign main_genericstandalone_rx_last_be_source_stb = main_genericstandalone_rx_last_be_sink_stb;
assign main_genericstandalone_rx_last_be_sink_ack = main_genericstandalone_rx_last_be_source_ack;
assign main_genericstandalone_rx_last_be_source_last = main_genericstandalone_rx_last_be_sink_last;
assign main_genericstandalone_rx_last_be_source_eop = main_genericstandalone_rx_last_be_sink_eop;
assign main_genericstandalone_rx_last_be_source_payload_data = main_genericstandalone_rx_last_be_sink_payload_data;
assign main_genericstandalone_rx_last_be_source_payload_error = main_genericstandalone_rx_last_be_sink_payload_error;

// synthesis translate_off
reg dummy_d_49;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_last_be_source_payload_last_be <= 1'd0;
	main_genericstandalone_rx_last_be_source_payload_last_be <= main_genericstandalone_rx_last_be_sink_payload_last_be;
	main_genericstandalone_rx_last_be_source_payload_last_be <= main_genericstandalone_rx_last_be_sink_eop;
// synthesis translate_off
	dummy_d_49 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_tx_converter_converter_sink_stb = main_genericstandalone_tx_converter_sink_sink_stb;
assign main_genericstandalone_tx_converter_converter_sink_last = main_genericstandalone_tx_converter_sink_sink_last;
assign main_genericstandalone_tx_converter_converter_sink_eop = main_genericstandalone_tx_converter_sink_sink_eop;
assign main_genericstandalone_tx_converter_sink_sink_ack = main_genericstandalone_tx_converter_converter_sink_ack;

// synthesis translate_off
reg dummy_d_50;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_converter_converter_sink_payload_data <= 80'd0;
	main_genericstandalone_tx_converter_converter_sink_payload_data[7:0] <= main_genericstandalone_tx_converter_sink_sink_payload_data[7:0];
	main_genericstandalone_tx_converter_converter_sink_payload_data[8] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[0];
	main_genericstandalone_tx_converter_converter_sink_payload_data[9] <= main_genericstandalone_tx_converter_sink_sink_payload_error[0];
	main_genericstandalone_tx_converter_converter_sink_payload_data[17:10] <= main_genericstandalone_tx_converter_sink_sink_payload_data[15:8];
	main_genericstandalone_tx_converter_converter_sink_payload_data[18] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[1];
	main_genericstandalone_tx_converter_converter_sink_payload_data[19] <= main_genericstandalone_tx_converter_sink_sink_payload_error[1];
	main_genericstandalone_tx_converter_converter_sink_payload_data[27:20] <= main_genericstandalone_tx_converter_sink_sink_payload_data[23:16];
	main_genericstandalone_tx_converter_converter_sink_payload_data[28] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[2];
	main_genericstandalone_tx_converter_converter_sink_payload_data[29] <= main_genericstandalone_tx_converter_sink_sink_payload_error[2];
	main_genericstandalone_tx_converter_converter_sink_payload_data[37:30] <= main_genericstandalone_tx_converter_sink_sink_payload_data[31:24];
	main_genericstandalone_tx_converter_converter_sink_payload_data[38] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[3];
	main_genericstandalone_tx_converter_converter_sink_payload_data[39] <= main_genericstandalone_tx_converter_sink_sink_payload_error[3];
	main_genericstandalone_tx_converter_converter_sink_payload_data[47:40] <= main_genericstandalone_tx_converter_sink_sink_payload_data[39:32];
	main_genericstandalone_tx_converter_converter_sink_payload_data[48] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[4];
	main_genericstandalone_tx_converter_converter_sink_payload_data[49] <= main_genericstandalone_tx_converter_sink_sink_payload_error[4];
	main_genericstandalone_tx_converter_converter_sink_payload_data[57:50] <= main_genericstandalone_tx_converter_sink_sink_payload_data[47:40];
	main_genericstandalone_tx_converter_converter_sink_payload_data[58] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[5];
	main_genericstandalone_tx_converter_converter_sink_payload_data[59] <= main_genericstandalone_tx_converter_sink_sink_payload_error[5];
	main_genericstandalone_tx_converter_converter_sink_payload_data[67:60] <= main_genericstandalone_tx_converter_sink_sink_payload_data[55:48];
	main_genericstandalone_tx_converter_converter_sink_payload_data[68] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[6];
	main_genericstandalone_tx_converter_converter_sink_payload_data[69] <= main_genericstandalone_tx_converter_sink_sink_payload_error[6];
	main_genericstandalone_tx_converter_converter_sink_payload_data[77:70] <= main_genericstandalone_tx_converter_sink_sink_payload_data[63:56];
	main_genericstandalone_tx_converter_converter_sink_payload_data[78] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[7];
	main_genericstandalone_tx_converter_converter_sink_payload_data[79] <= main_genericstandalone_tx_converter_sink_sink_payload_error[7];
// synthesis translate_off
	dummy_d_50 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_tx_converter_source_source_stb = main_genericstandalone_tx_converter_converter_source_stb;
assign main_genericstandalone_tx_converter_source_source_last = main_genericstandalone_tx_converter_converter_source_last;
assign main_genericstandalone_tx_converter_source_source_eop = main_genericstandalone_tx_converter_converter_source_eop;
assign main_genericstandalone_tx_converter_converter_source_ack = main_genericstandalone_tx_converter_source_source_ack;
assign {main_genericstandalone_tx_converter_source_source_payload_error, main_genericstandalone_tx_converter_source_source_payload_last_be, main_genericstandalone_tx_converter_source_source_payload_data} = main_genericstandalone_tx_converter_converter_source_payload_data;
assign main_genericstandalone_tx_converter_converter_last = (main_genericstandalone_tx_converter_converter_mux == 3'd7);
assign main_genericstandalone_tx_converter_converter_source_stb = main_genericstandalone_tx_converter_converter_sink_stb;
assign main_genericstandalone_tx_converter_converter_source_eop = (main_genericstandalone_tx_converter_converter_sink_eop & main_genericstandalone_tx_converter_converter_last);
assign main_genericstandalone_tx_converter_converter_source_last = (main_genericstandalone_tx_converter_converter_sink_last & main_genericstandalone_tx_converter_converter_last);
assign main_genericstandalone_tx_converter_converter_sink_ack = (main_genericstandalone_tx_converter_converter_last & main_genericstandalone_tx_converter_converter_source_ack);

// synthesis translate_off
reg dummy_d_51;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_converter_converter_source_payload_data <= 10'd0;
	case (main_genericstandalone_tx_converter_converter_mux)
		1'd0: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[9:0];
		end
		1'd1: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[19:10];
		end
		2'd2: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[29:20];
		end
		2'd3: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[39:30];
		end
		3'd4: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[49:40];
		end
		3'd5: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[59:50];
		end
		3'd6: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[69:60];
		end
		default: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[79:70];
		end
	endcase
// synthesis translate_off
	dummy_d_51 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_converter_converter_sink_stb = main_genericstandalone_rx_converter_sink_sink_stb;
assign main_genericstandalone_rx_converter_converter_sink_last = main_genericstandalone_rx_converter_sink_sink_last;
assign main_genericstandalone_rx_converter_converter_sink_eop = main_genericstandalone_rx_converter_sink_sink_eop;
assign main_genericstandalone_rx_converter_sink_sink_ack = main_genericstandalone_rx_converter_converter_sink_ack;
assign main_genericstandalone_rx_converter_converter_sink_payload_data = {main_genericstandalone_rx_converter_sink_sink_payload_error, main_genericstandalone_rx_converter_sink_sink_payload_last_be, main_genericstandalone_rx_converter_sink_sink_payload_data};
assign main_genericstandalone_rx_converter_source_source_stb = main_genericstandalone_rx_converter_converter_source_stb;
assign main_genericstandalone_rx_converter_source_source_last = main_genericstandalone_rx_converter_converter_source_last;
assign main_genericstandalone_rx_converter_source_source_eop = main_genericstandalone_rx_converter_converter_source_eop;
assign main_genericstandalone_rx_converter_converter_source_ack = main_genericstandalone_rx_converter_source_source_ack;

// synthesis translate_off
reg dummy_d_52;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_converter_source_source_payload_data <= 64'd0;
	main_genericstandalone_rx_converter_source_source_payload_data[7:0] <= main_genericstandalone_rx_converter_converter_source_payload_data[7:0];
	main_genericstandalone_rx_converter_source_source_payload_data[15:8] <= main_genericstandalone_rx_converter_converter_source_payload_data[17:10];
	main_genericstandalone_rx_converter_source_source_payload_data[23:16] <= main_genericstandalone_rx_converter_converter_source_payload_data[27:20];
	main_genericstandalone_rx_converter_source_source_payload_data[31:24] <= main_genericstandalone_rx_converter_converter_source_payload_data[37:30];
	main_genericstandalone_rx_converter_source_source_payload_data[39:32] <= main_genericstandalone_rx_converter_converter_source_payload_data[47:40];
	main_genericstandalone_rx_converter_source_source_payload_data[47:40] <= main_genericstandalone_rx_converter_converter_source_payload_data[57:50];
	main_genericstandalone_rx_converter_source_source_payload_data[55:48] <= main_genericstandalone_rx_converter_converter_source_payload_data[67:60];
	main_genericstandalone_rx_converter_source_source_payload_data[63:56] <= main_genericstandalone_rx_converter_converter_source_payload_data[77:70];
// synthesis translate_off
	dummy_d_52 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_53;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_converter_source_source_payload_last_be <= 8'd0;
	main_genericstandalone_rx_converter_source_source_payload_last_be[0] <= main_genericstandalone_rx_converter_converter_source_payload_data[8];
	main_genericstandalone_rx_converter_source_source_payload_last_be[1] <= main_genericstandalone_rx_converter_converter_source_payload_data[18];
	main_genericstandalone_rx_converter_source_source_payload_last_be[2] <= main_genericstandalone_rx_converter_converter_source_payload_data[28];
	main_genericstandalone_rx_converter_source_source_payload_last_be[3] <= main_genericstandalone_rx_converter_converter_source_payload_data[38];
	main_genericstandalone_rx_converter_source_source_payload_last_be[4] <= main_genericstandalone_rx_converter_converter_source_payload_data[48];
	main_genericstandalone_rx_converter_source_source_payload_last_be[5] <= main_genericstandalone_rx_converter_converter_source_payload_data[58];
	main_genericstandalone_rx_converter_source_source_payload_last_be[6] <= main_genericstandalone_rx_converter_converter_source_payload_data[68];
	main_genericstandalone_rx_converter_source_source_payload_last_be[7] <= main_genericstandalone_rx_converter_converter_source_payload_data[78];
// synthesis translate_off
	dummy_d_53 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_54;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_converter_source_source_payload_error <= 8'd0;
	main_genericstandalone_rx_converter_source_source_payload_error[0] <= main_genericstandalone_rx_converter_converter_source_payload_data[9];
	main_genericstandalone_rx_converter_source_source_payload_error[1] <= main_genericstandalone_rx_converter_converter_source_payload_data[19];
	main_genericstandalone_rx_converter_source_source_payload_error[2] <= main_genericstandalone_rx_converter_converter_source_payload_data[29];
	main_genericstandalone_rx_converter_source_source_payload_error[3] <= main_genericstandalone_rx_converter_converter_source_payload_data[39];
	main_genericstandalone_rx_converter_source_source_payload_error[4] <= main_genericstandalone_rx_converter_converter_source_payload_data[49];
	main_genericstandalone_rx_converter_source_source_payload_error[5] <= main_genericstandalone_rx_converter_converter_source_payload_data[59];
	main_genericstandalone_rx_converter_source_source_payload_error[6] <= main_genericstandalone_rx_converter_converter_source_payload_data[69];
	main_genericstandalone_rx_converter_source_source_payload_error[7] <= main_genericstandalone_rx_converter_converter_source_payload_data[79];
// synthesis translate_off
	dummy_d_54 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_converter_converter_sink_ack = ((~main_genericstandalone_rx_converter_converter_strobe_all) | main_genericstandalone_rx_converter_converter_source_ack);
assign main_genericstandalone_rx_converter_converter_source_stb = main_genericstandalone_rx_converter_converter_strobe_all;
assign main_genericstandalone_rx_converter_converter_load_part = (main_genericstandalone_rx_converter_converter_sink_stb & main_genericstandalone_rx_converter_converter_sink_ack);
assign main_genericstandalone_rx_converter_converter_source_last = 1'd1;
assign main_genericstandalone_tx_cdc_asyncfifo_din = {main_genericstandalone_tx_cdc_fifo_in_eop, main_genericstandalone_tx_cdc_fifo_in_payload_error, main_genericstandalone_tx_cdc_fifo_in_payload_last_be, main_genericstandalone_tx_cdc_fifo_in_payload_data};
assign {main_genericstandalone_tx_cdc_fifo_out_eop, main_genericstandalone_tx_cdc_fifo_out_payload_error, main_genericstandalone_tx_cdc_fifo_out_payload_last_be, main_genericstandalone_tx_cdc_fifo_out_payload_data} = main_genericstandalone_tx_cdc_asyncfifo_dout;
assign main_genericstandalone_tx_cdc_sink_ack = main_genericstandalone_tx_cdc_asyncfifo_writable;
assign main_genericstandalone_tx_cdc_asyncfifo_we = main_genericstandalone_tx_cdc_sink_stb;
assign main_genericstandalone_tx_cdc_fifo_in_eop = main_genericstandalone_tx_cdc_sink_eop;
assign main_genericstandalone_tx_cdc_fifo_in_payload_data = main_genericstandalone_tx_cdc_sink_payload_data;
assign main_genericstandalone_tx_cdc_fifo_in_payload_last_be = main_genericstandalone_tx_cdc_sink_payload_last_be;
assign main_genericstandalone_tx_cdc_fifo_in_payload_error = main_genericstandalone_tx_cdc_sink_payload_error;
assign main_genericstandalone_tx_cdc_source_stb = main_genericstandalone_tx_cdc_asyncfifo_readable;
assign main_genericstandalone_tx_cdc_source_eop = main_genericstandalone_tx_cdc_fifo_out_eop;
assign main_genericstandalone_tx_cdc_source_payload_data = main_genericstandalone_tx_cdc_fifo_out_payload_data;
assign main_genericstandalone_tx_cdc_source_payload_last_be = main_genericstandalone_tx_cdc_fifo_out_payload_last_be;
assign main_genericstandalone_tx_cdc_source_payload_error = main_genericstandalone_tx_cdc_fifo_out_payload_error;
assign main_genericstandalone_tx_cdc_asyncfifo_re = main_genericstandalone_tx_cdc_source_ack;
assign main_genericstandalone_tx_cdc_graycounter0_ce = (main_genericstandalone_tx_cdc_asyncfifo_writable & main_genericstandalone_tx_cdc_asyncfifo_we);
assign main_genericstandalone_tx_cdc_graycounter1_ce = (main_genericstandalone_tx_cdc_asyncfifo_readable & main_genericstandalone_tx_cdc_asyncfifo_re);
assign main_genericstandalone_tx_cdc_asyncfifo_writable = (((main_genericstandalone_tx_cdc_graycounter0_q[6] == main_genericstandalone_tx_cdc_consume_wdomain[6]) | (main_genericstandalone_tx_cdc_graycounter0_q[5] == main_genericstandalone_tx_cdc_consume_wdomain[5])) | (main_genericstandalone_tx_cdc_graycounter0_q[4:0] != main_genericstandalone_tx_cdc_consume_wdomain[4:0]));
assign main_genericstandalone_tx_cdc_asyncfifo_readable = (main_genericstandalone_tx_cdc_graycounter1_q != main_genericstandalone_tx_cdc_produce_rdomain);
assign main_genericstandalone_tx_cdc_wrport_adr = main_genericstandalone_tx_cdc_graycounter0_q_binary[5:0];
assign main_genericstandalone_tx_cdc_wrport_dat_w = main_genericstandalone_tx_cdc_asyncfifo_din;
assign main_genericstandalone_tx_cdc_wrport_we = main_genericstandalone_tx_cdc_graycounter0_ce;
assign main_genericstandalone_tx_cdc_rdport_adr = main_genericstandalone_tx_cdc_graycounter1_q_next_binary[5:0];
assign main_genericstandalone_tx_cdc_asyncfifo_dout = main_genericstandalone_tx_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_55;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (main_genericstandalone_tx_cdc_graycounter0_ce) begin
		main_genericstandalone_tx_cdc_graycounter0_q_next_binary <= (main_genericstandalone_tx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		main_genericstandalone_tx_cdc_graycounter0_q_next_binary <= main_genericstandalone_tx_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_55 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_tx_cdc_graycounter0_q_next = (main_genericstandalone_tx_cdc_graycounter0_q_next_binary ^ main_genericstandalone_tx_cdc_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_56;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (main_genericstandalone_tx_cdc_graycounter1_ce) begin
		main_genericstandalone_tx_cdc_graycounter1_q_next_binary <= (main_genericstandalone_tx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		main_genericstandalone_tx_cdc_graycounter1_q_next_binary <= main_genericstandalone_tx_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_56 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_tx_cdc_graycounter1_q_next = (main_genericstandalone_tx_cdc_graycounter1_q_next_binary ^ main_genericstandalone_tx_cdc_graycounter1_q_next_binary[6:1]);
assign main_genericstandalone_rx_cdc_asyncfifo_din = {main_genericstandalone_rx_cdc_fifo_in_eop, main_genericstandalone_rx_cdc_fifo_in_payload_error, main_genericstandalone_rx_cdc_fifo_in_payload_last_be, main_genericstandalone_rx_cdc_fifo_in_payload_data};
assign {main_genericstandalone_rx_cdc_fifo_out_eop, main_genericstandalone_rx_cdc_fifo_out_payload_error, main_genericstandalone_rx_cdc_fifo_out_payload_last_be, main_genericstandalone_rx_cdc_fifo_out_payload_data} = main_genericstandalone_rx_cdc_asyncfifo_dout;
assign main_genericstandalone_rx_cdc_sink_ack = main_genericstandalone_rx_cdc_asyncfifo_writable;
assign main_genericstandalone_rx_cdc_asyncfifo_we = main_genericstandalone_rx_cdc_sink_stb;
assign main_genericstandalone_rx_cdc_fifo_in_eop = main_genericstandalone_rx_cdc_sink_eop;
assign main_genericstandalone_rx_cdc_fifo_in_payload_data = main_genericstandalone_rx_cdc_sink_payload_data;
assign main_genericstandalone_rx_cdc_fifo_in_payload_last_be = main_genericstandalone_rx_cdc_sink_payload_last_be;
assign main_genericstandalone_rx_cdc_fifo_in_payload_error = main_genericstandalone_rx_cdc_sink_payload_error;
assign main_genericstandalone_rx_cdc_source_stb = main_genericstandalone_rx_cdc_asyncfifo_readable;
assign main_genericstandalone_rx_cdc_source_eop = main_genericstandalone_rx_cdc_fifo_out_eop;
assign main_genericstandalone_rx_cdc_source_payload_data = main_genericstandalone_rx_cdc_fifo_out_payload_data;
assign main_genericstandalone_rx_cdc_source_payload_last_be = main_genericstandalone_rx_cdc_fifo_out_payload_last_be;
assign main_genericstandalone_rx_cdc_source_payload_error = main_genericstandalone_rx_cdc_fifo_out_payload_error;
assign main_genericstandalone_rx_cdc_asyncfifo_re = main_genericstandalone_rx_cdc_source_ack;
assign main_genericstandalone_rx_cdc_graycounter0_ce = (main_genericstandalone_rx_cdc_asyncfifo_writable & main_genericstandalone_rx_cdc_asyncfifo_we);
assign main_genericstandalone_rx_cdc_graycounter1_ce = (main_genericstandalone_rx_cdc_asyncfifo_readable & main_genericstandalone_rx_cdc_asyncfifo_re);
assign main_genericstandalone_rx_cdc_asyncfifo_writable = (((main_genericstandalone_rx_cdc_graycounter0_q[6] == main_genericstandalone_rx_cdc_consume_wdomain[6]) | (main_genericstandalone_rx_cdc_graycounter0_q[5] == main_genericstandalone_rx_cdc_consume_wdomain[5])) | (main_genericstandalone_rx_cdc_graycounter0_q[4:0] != main_genericstandalone_rx_cdc_consume_wdomain[4:0]));
assign main_genericstandalone_rx_cdc_asyncfifo_readable = (main_genericstandalone_rx_cdc_graycounter1_q != main_genericstandalone_rx_cdc_produce_rdomain);
assign main_genericstandalone_rx_cdc_wrport_adr = main_genericstandalone_rx_cdc_graycounter0_q_binary[5:0];
assign main_genericstandalone_rx_cdc_wrport_dat_w = main_genericstandalone_rx_cdc_asyncfifo_din;
assign main_genericstandalone_rx_cdc_wrport_we = main_genericstandalone_rx_cdc_graycounter0_ce;
assign main_genericstandalone_rx_cdc_rdport_adr = main_genericstandalone_rx_cdc_graycounter1_q_next_binary[5:0];
assign main_genericstandalone_rx_cdc_asyncfifo_dout = main_genericstandalone_rx_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_57;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (main_genericstandalone_rx_cdc_graycounter0_ce) begin
		main_genericstandalone_rx_cdc_graycounter0_q_next_binary <= (main_genericstandalone_rx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		main_genericstandalone_rx_cdc_graycounter0_q_next_binary <= main_genericstandalone_rx_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_57 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_cdc_graycounter0_q_next = (main_genericstandalone_rx_cdc_graycounter0_q_next_binary ^ main_genericstandalone_rx_cdc_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_58;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (main_genericstandalone_rx_cdc_graycounter1_ce) begin
		main_genericstandalone_rx_cdc_graycounter1_q_next_binary <= (main_genericstandalone_rx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		main_genericstandalone_rx_cdc_graycounter1_q_next_binary <= main_genericstandalone_rx_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_58 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_cdc_graycounter1_q_next = (main_genericstandalone_rx_cdc_graycounter1_q_next_binary ^ main_genericstandalone_rx_cdc_graycounter1_q_next_binary[6:1]);
assign main_genericstandalone_sram8_sink_stb = main_genericstandalone_sink_sink_stb;
assign main_genericstandalone_sink_sink_ack = main_genericstandalone_sram9_sink_ack;
assign main_genericstandalone_sram10_sink_last = main_genericstandalone_sink_sink_last;
assign main_genericstandalone_sram11_sink_eop = main_genericstandalone_sink_sink_eop;
assign main_genericstandalone_sram12_sink_payload_data = main_genericstandalone_sink_sink_payload_data;
assign main_genericstandalone_sram13_sink_payload_last_be = main_genericstandalone_sink_sink_payload_last_be;
assign main_genericstandalone_sram14_sink_payload_error = main_genericstandalone_sink_sink_payload_error;
assign main_genericstandalone_source_source_stb = main_genericstandalone_sram88_source_stb;
assign main_genericstandalone_sram89_source_ack = main_genericstandalone_source_source_ack;
assign main_genericstandalone_source_source_last = main_genericstandalone_sram90_source_last;
assign main_genericstandalone_source_source_eop = main_genericstandalone_sram91_source_eop;
assign main_genericstandalone_source_source_payload_data = main_genericstandalone_sram92_source_payload_data;
assign main_genericstandalone_source_source_payload_last_be = main_genericstandalone_sram93_source_payload_last_be;
assign main_genericstandalone_source_source_payload_error = main_genericstandalone_sram94_source_payload_error;
assign main_genericstandalone_sram42_sink_payload_slot = main_genericstandalone_slot;
assign main_genericstandalone_sram43_sink_payload_length = main_genericstandalone_sram33_counter;
assign main_genericstandalone_sram45_source_ack = main_genericstandalone_sram22_clear;
assign main_genericstandalone_sram21_trigger = main_genericstandalone_sram44_source_stb;
assign main_genericstandalone_sram15_status = main_genericstandalone_sram47_source_payload_slot;
assign main_genericstandalone_sram16_status = main_genericstandalone_sram48_source_payload_length;

// synthesis translate_off
reg dummy_d_59;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram72_adr <= 8'd0;
	main_genericstandalone_sram74_we <= 1'd0;
	main_genericstandalone_sram75_dat_w <= 64'd0;
	main_genericstandalone_sram76_adr <= 8'd0;
	main_genericstandalone_sram78_we <= 1'd0;
	main_genericstandalone_sram79_dat_w <= 64'd0;
	main_genericstandalone_sram80_adr <= 8'd0;
	main_genericstandalone_sram82_we <= 1'd0;
	main_genericstandalone_sram83_dat_w <= 64'd0;
	main_genericstandalone_sram84_adr <= 8'd0;
	main_genericstandalone_sram86_we <= 1'd0;
	main_genericstandalone_sram87_dat_w <= 64'd0;
	case (main_genericstandalone_slot)
		1'd0: begin
			main_genericstandalone_sram72_adr <= main_genericstandalone_sram33_counter[10:3];
			main_genericstandalone_sram75_dat_w <= main_genericstandalone_sram12_sink_payload_data;
			if ((main_genericstandalone_sram8_sink_stb & main_genericstandalone_ongoing)) begin
				main_genericstandalone_sram74_we <= 4'd15;
			end
		end
		1'd1: begin
			main_genericstandalone_sram76_adr <= main_genericstandalone_sram33_counter[10:3];
			main_genericstandalone_sram79_dat_w <= main_genericstandalone_sram12_sink_payload_data;
			if ((main_genericstandalone_sram8_sink_stb & main_genericstandalone_ongoing)) begin
				main_genericstandalone_sram78_we <= 4'd15;
			end
		end
		2'd2: begin
			main_genericstandalone_sram80_adr <= main_genericstandalone_sram33_counter[10:3];
			main_genericstandalone_sram83_dat_w <= main_genericstandalone_sram12_sink_payload_data;
			if ((main_genericstandalone_sram8_sink_stb & main_genericstandalone_ongoing)) begin
				main_genericstandalone_sram82_we <= 4'd15;
			end
		end
		2'd3: begin
			main_genericstandalone_sram84_adr <= main_genericstandalone_sram33_counter[10:3];
			main_genericstandalone_sram87_dat_w <= main_genericstandalone_sram12_sink_payload_data;
			if ((main_genericstandalone_sram8_sink_stb & main_genericstandalone_ongoing)) begin
				main_genericstandalone_sram86_we <= 4'd15;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_59 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram25_status_w = main_genericstandalone_sram19_status;

// synthesis translate_off
reg dummy_d_60;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram22_clear <= 1'd0;
	if ((main_genericstandalone_sram26_pending_re & main_genericstandalone_sram27_pending_r)) begin
		main_genericstandalone_sram22_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_60 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram28_pending_w = main_genericstandalone_sram20_pending;
assign main_genericstandalone_sram18_irq = (main_genericstandalone_sram28_pending_w & main_genericstandalone_sram30_storage);
assign main_genericstandalone_sram19_status = main_genericstandalone_sram21_trigger;
assign main_genericstandalone_sram20_pending = main_genericstandalone_sram21_trigger;

// synthesis translate_off
reg dummy_d_61;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_decoded <= 4'd0;
	case (main_genericstandalone_sram13_sink_payload_last_be)
		1'd1: begin
			main_genericstandalone_decoded <= 1'd1;
		end
		2'd2: begin
			main_genericstandalone_decoded <= 2'd2;
		end
		3'd4: begin
			main_genericstandalone_decoded <= 2'd3;
		end
		4'd8: begin
			main_genericstandalone_decoded <= 3'd4;
		end
		5'd16: begin
			main_genericstandalone_decoded <= 3'd5;
		end
		6'd32: begin
			main_genericstandalone_decoded <= 3'd6;
		end
		7'd64: begin
			main_genericstandalone_decoded <= 3'd7;
		end
		default: begin
			main_genericstandalone_decoded <= 4'd8;
		end
	endcase
// synthesis translate_off
	dummy_d_61 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram53_din = {main_genericstandalone_sram68_fifo_in_eop, main_genericstandalone_sram67_fifo_in_payload_length, main_genericstandalone_sram66_fifo_in_payload_slot};
assign {main_genericstandalone_sram71_fifo_out_eop, main_genericstandalone_sram70_fifo_out_payload_length, main_genericstandalone_sram69_fifo_out_payload_slot} = main_genericstandalone_sram54_dout;
assign main_genericstandalone_sram40_sink_ack = main_genericstandalone_sram50_writable;
assign main_genericstandalone_sram49_we = main_genericstandalone_sram39_sink_stb;
assign main_genericstandalone_sram68_fifo_in_eop = main_genericstandalone_sram41_sink_eop;
assign main_genericstandalone_sram66_fifo_in_payload_slot = main_genericstandalone_sram42_sink_payload_slot;
assign main_genericstandalone_sram67_fifo_in_payload_length = main_genericstandalone_sram43_sink_payload_length;
assign main_genericstandalone_sram44_source_stb = main_genericstandalone_sram52_readable;
assign main_genericstandalone_sram46_source_eop = main_genericstandalone_sram71_fifo_out_eop;
assign main_genericstandalone_sram47_source_payload_slot = main_genericstandalone_sram69_fifo_out_payload_slot;
assign main_genericstandalone_sram48_source_payload_length = main_genericstandalone_sram70_fifo_out_payload_length;
assign main_genericstandalone_sram51_re = main_genericstandalone_sram45_source_ack;

// synthesis translate_off
reg dummy_d_62;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram59_adr <= 2'd0;
	if (main_genericstandalone_sram56_replace) begin
		main_genericstandalone_sram59_adr <= (main_genericstandalone_sram57_produce - 1'd1);
	end else begin
		main_genericstandalone_sram59_adr <= main_genericstandalone_sram57_produce;
	end
// synthesis translate_off
	dummy_d_62 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram62_dat_w = main_genericstandalone_sram53_din;
assign main_genericstandalone_sram61_we = (main_genericstandalone_sram49_we & (main_genericstandalone_sram50_writable | main_genericstandalone_sram56_replace));
assign main_genericstandalone_sram63_do_read = (main_genericstandalone_sram52_readable & main_genericstandalone_sram51_re);
assign main_genericstandalone_sram64_adr = main_genericstandalone_sram58_consume;
assign main_genericstandalone_sram54_dout = main_genericstandalone_sram65_dat_r;
assign main_genericstandalone_sram50_writable = (main_genericstandalone_sram55_level != 3'd4);
assign main_genericstandalone_sram52_readable = (main_genericstandalone_sram55_level != 1'd0);

// synthesis translate_off
reg dummy_d_63;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram34_counter_reset <= 1'd0;
	main_genericstandalone_sram35_counter_ce <= 1'd0;
	main_genericstandalone_slot_ce <= 1'd0;
	main_genericstandalone_ongoing <= 1'd0;
	main_genericstandalone_sram39_sink_stb <= 1'd0;
	builder_liteethmacsramwriter_next_state <= 2'd0;
	main_genericstandalone_sram17_status_liteethmac_next_value <= 32'd0;
	main_genericstandalone_sram17_status_liteethmac_next_value_ce <= 1'd0;
	builder_liteethmacsramwriter_next_state <= builder_liteethmacsramwriter_state;
	case (builder_liteethmacsramwriter_state)
		1'd1: begin
			if (main_genericstandalone_sram8_sink_stb) begin
				if ((main_genericstandalone_sram33_counter == 11'd1530)) begin
					builder_liteethmacsramwriter_next_state <= 2'd2;
				end else begin
					main_genericstandalone_sram35_counter_ce <= 1'd1;
					main_genericstandalone_ongoing <= 1'd1;
				end
				if (main_genericstandalone_sram11_sink_eop) begin
					if (((main_genericstandalone_sram14_sink_payload_error & main_genericstandalone_sram13_sink_payload_last_be) != 1'd0)) begin
						main_genericstandalone_sram34_counter_reset <= 1'd1;
						builder_liteethmacsramwriter_next_state <= 1'd0;
					end else begin
						builder_liteethmacsramwriter_next_state <= 2'd3;
					end
				end
			end
		end
		2'd2: begin
			main_genericstandalone_sram34_counter_reset <= 1'd1;
			if ((main_genericstandalone_sram8_sink_stb & main_genericstandalone_sram11_sink_eop)) begin
				main_genericstandalone_sram17_status_liteethmac_next_value <= (main_genericstandalone_sram17_status + 1'd1);
				main_genericstandalone_sram17_status_liteethmac_next_value_ce <= 1'd1;
				builder_liteethmacsramwriter_next_state <= 1'd0;
			end
		end
		2'd3: begin
			main_genericstandalone_sram34_counter_reset <= 1'd1;
			main_genericstandalone_slot_ce <= 1'd1;
			main_genericstandalone_sram39_sink_stb <= 1'd1;
			builder_liteethmacsramwriter_next_state <= 1'd0;
		end
		default: begin
			if (main_genericstandalone_sram8_sink_stb) begin
				if (main_genericstandalone_sram40_sink_ack) begin
					main_genericstandalone_ongoing <= 1'd1;
					main_genericstandalone_sram35_counter_ce <= 1'd1;
					builder_liteethmacsramwriter_next_state <= 1'd1;
				end else begin
					builder_liteethmacsramwriter_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_63 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram119_sink_stb = main_genericstandalone_start_re;
assign main_genericstandalone_sram122_sink_payload_slot = main_genericstandalone_sram100_storage;
assign main_genericstandalone_sram123_sink_payload_length = main_genericstandalone_sram103_storage;
assign main_genericstandalone_sram98_status = main_genericstandalone_sram120_sink_ack;

// synthesis translate_off
reg dummy_d_64;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram93_source_payload_last_be <= 8'd0;
	if (main_genericstandalone_last) begin
		main_genericstandalone_sram93_source_payload_last_be <= main_genericstandalone_encoded;
	end
// synthesis translate_off
	dummy_d_64 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_last = ((main_genericstandalone_sram152_counter + 4'd8) >= main_genericstandalone_sram128_source_payload_length);
assign main_genericstandalone_sram158_adr = main_genericstandalone_sram152_counter[10:3];
assign main_genericstandalone_sram160_adr = main_genericstandalone_sram152_counter[10:3];
assign main_genericstandalone_sram162_adr = main_genericstandalone_sram152_counter[10:3];
assign main_genericstandalone_sram164_adr = main_genericstandalone_sram152_counter[10:3];

// synthesis translate_off
reg dummy_d_65;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram92_source_payload_data <= 64'd0;
	case (main_genericstandalone_sram127_source_payload_slot)
		1'd0: begin
			main_genericstandalone_sram92_source_payload_data <= main_genericstandalone_sram159_dat_r;
		end
		1'd1: begin
			main_genericstandalone_sram92_source_payload_data <= main_genericstandalone_sram161_dat_r;
		end
		2'd2: begin
			main_genericstandalone_sram92_source_payload_data <= main_genericstandalone_sram163_dat_r;
		end
		2'd3: begin
			main_genericstandalone_sram92_source_payload_data <= main_genericstandalone_sram165_dat_r;
		end
	endcase
// synthesis translate_off
	dummy_d_65 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram112_status_w = main_genericstandalone_sram106_status;

// synthesis translate_off
reg dummy_d_66;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram109_clear <= 1'd0;
	if ((main_genericstandalone_sram113_pending_re & main_genericstandalone_sram114_pending_r)) begin
		main_genericstandalone_sram109_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_66 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram115_pending_w = main_genericstandalone_sram107_pending;
assign main_genericstandalone_sram105_irq = (main_genericstandalone_sram115_pending_w & main_genericstandalone_sram117_storage);
assign main_genericstandalone_sram106_status = 1'd0;
assign main_genericstandalone_sram133_din = {main_genericstandalone_sram148_fifo_in_eop, main_genericstandalone_sram147_fifo_in_payload_length, main_genericstandalone_sram146_fifo_in_payload_slot};
assign {main_genericstandalone_sram151_fifo_out_eop, main_genericstandalone_sram150_fifo_out_payload_length, main_genericstandalone_sram149_fifo_out_payload_slot} = main_genericstandalone_sram134_dout;
assign main_genericstandalone_sram120_sink_ack = main_genericstandalone_sram130_writable;
assign main_genericstandalone_sram129_we = main_genericstandalone_sram119_sink_stb;
assign main_genericstandalone_sram148_fifo_in_eop = main_genericstandalone_sram121_sink_eop;
assign main_genericstandalone_sram146_fifo_in_payload_slot = main_genericstandalone_sram122_sink_payload_slot;
assign main_genericstandalone_sram147_fifo_in_payload_length = main_genericstandalone_sram123_sink_payload_length;
assign main_genericstandalone_sram124_source_stb = main_genericstandalone_sram132_readable;
assign main_genericstandalone_sram126_source_eop = main_genericstandalone_sram151_fifo_out_eop;
assign main_genericstandalone_sram127_source_payload_slot = main_genericstandalone_sram149_fifo_out_payload_slot;
assign main_genericstandalone_sram128_source_payload_length = main_genericstandalone_sram150_fifo_out_payload_length;
assign main_genericstandalone_sram131_re = main_genericstandalone_sram125_source_ack;

// synthesis translate_off
reg dummy_d_67;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram139_adr <= 2'd0;
	if (main_genericstandalone_sram136_replace) begin
		main_genericstandalone_sram139_adr <= (main_genericstandalone_sram137_produce - 1'd1);
	end else begin
		main_genericstandalone_sram139_adr <= main_genericstandalone_sram137_produce;
	end
// synthesis translate_off
	dummy_d_67 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram142_dat_w = main_genericstandalone_sram133_din;
assign main_genericstandalone_sram141_we = (main_genericstandalone_sram129_we & (main_genericstandalone_sram130_writable | main_genericstandalone_sram136_replace));
assign main_genericstandalone_sram143_do_read = (main_genericstandalone_sram132_readable & main_genericstandalone_sram131_re);
assign main_genericstandalone_sram144_adr = main_genericstandalone_sram138_consume;
assign main_genericstandalone_sram134_dout = main_genericstandalone_sram145_dat_r;
assign main_genericstandalone_sram130_writable = (main_genericstandalone_sram135_level != 3'd4);
assign main_genericstandalone_sram132_readable = (main_genericstandalone_sram135_level != 1'd0);

// synthesis translate_off
reg dummy_d_68;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram88_source_stb <= 1'd0;
	main_genericstandalone_sram91_source_eop <= 1'd0;
	main_genericstandalone_sram108_trigger <= 1'd0;
	main_genericstandalone_sram125_source_ack <= 1'd0;
	main_genericstandalone_sram153_counter_reset <= 1'd0;
	main_genericstandalone_sram154_counter_ce <= 1'd0;
	builder_liteethmacsramreader_next_state <= 2'd0;
	builder_liteethmacsramreader_next_state <= builder_liteethmacsramreader_state;
	case (builder_liteethmacsramreader_state)
		1'd1: begin
			if ((~main_genericstandalone_last_d)) begin
				builder_liteethmacsramreader_next_state <= 2'd2;
			end else begin
				builder_liteethmacsramreader_next_state <= 2'd3;
			end
		end
		2'd2: begin
			main_genericstandalone_sram88_source_stb <= 1'd1;
			main_genericstandalone_sram91_source_eop <= main_genericstandalone_last;
			if (main_genericstandalone_sram89_source_ack) begin
				main_genericstandalone_sram154_counter_ce <= (~main_genericstandalone_last);
				builder_liteethmacsramreader_next_state <= 1'd1;
			end
		end
		2'd3: begin
			main_genericstandalone_sram125_source_ack <= 1'd1;
			main_genericstandalone_sram108_trigger <= 1'd1;
			builder_liteethmacsramreader_next_state <= 1'd0;
		end
		default: begin
			main_genericstandalone_sram153_counter_reset <= 1'd1;
			if (main_genericstandalone_sram124_source_stb) begin
				builder_liteethmacsramreader_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_68 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_69;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_encoded <= 8'd0;
	case (main_genericstandalone_sram128_source_payload_length[2:0])
		1'd1: begin
			main_genericstandalone_encoded <= 1'd1;
		end
		2'd2: begin
			main_genericstandalone_encoded <= 2'd2;
		end
		2'd3: begin
			main_genericstandalone_encoded <= 3'd4;
		end
		3'd4: begin
			main_genericstandalone_encoded <= 4'd8;
		end
		3'd5: begin
			main_genericstandalone_encoded <= 5'd16;
		end
		3'd6: begin
			main_genericstandalone_encoded <= 6'd32;
		end
		3'd7: begin
			main_genericstandalone_encoded <= 7'd64;
		end
		default: begin
			main_genericstandalone_encoded <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_69 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram166_irq = (main_genericstandalone_sram18_irq | main_genericstandalone_sram105_irq);
assign main_genericstandalone_sram0_adr = main_genericstandalone_sram0_bus_adr[7:0];
assign main_genericstandalone_sram0_bus_dat_r = main_genericstandalone_sram0_dat_r;
assign main_genericstandalone_sram1_adr = main_genericstandalone_sram1_bus_adr[7:0];
assign main_genericstandalone_sram1_bus_dat_r = main_genericstandalone_sram1_dat_r;
assign main_genericstandalone_sram2_adr = main_genericstandalone_sram2_bus_adr[7:0];
assign main_genericstandalone_sram2_bus_dat_r = main_genericstandalone_sram2_dat_r;
assign main_genericstandalone_sram3_adr = main_genericstandalone_sram3_bus_adr[7:0];
assign main_genericstandalone_sram3_bus_dat_r = main_genericstandalone_sram3_dat_r;

// synthesis translate_off
reg dummy_d_70;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram4_we <= 8'd0;
	main_genericstandalone_sram4_we[0] <= (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & main_genericstandalone_sram4_bus_we) & main_genericstandalone_sram4_bus_sel[0]);
	main_genericstandalone_sram4_we[1] <= (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & main_genericstandalone_sram4_bus_we) & main_genericstandalone_sram4_bus_sel[1]);
	main_genericstandalone_sram4_we[2] <= (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & main_genericstandalone_sram4_bus_we) & main_genericstandalone_sram4_bus_sel[2]);
	main_genericstandalone_sram4_we[3] <= (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & main_genericstandalone_sram4_bus_we) & main_genericstandalone_sram4_bus_sel[3]);
	main_genericstandalone_sram4_we[4] <= (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & main_genericstandalone_sram4_bus_we) & main_genericstandalone_sram4_bus_sel[4]);
	main_genericstandalone_sram4_we[5] <= (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & main_genericstandalone_sram4_bus_we) & main_genericstandalone_sram4_bus_sel[5]);
	main_genericstandalone_sram4_we[6] <= (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & main_genericstandalone_sram4_bus_we) & main_genericstandalone_sram4_bus_sel[6]);
	main_genericstandalone_sram4_we[7] <= (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & main_genericstandalone_sram4_bus_we) & main_genericstandalone_sram4_bus_sel[7]);
// synthesis translate_off
	dummy_d_70 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram4_adr = main_genericstandalone_sram4_bus_adr[7:0];
assign main_genericstandalone_sram4_bus_dat_r = main_genericstandalone_sram4_dat_r;
assign main_genericstandalone_sram4_dat_w = main_genericstandalone_sram4_bus_dat_w;

// synthesis translate_off
reg dummy_d_71;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram5_we <= 8'd0;
	main_genericstandalone_sram5_we[0] <= (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & main_genericstandalone_sram5_bus_we) & main_genericstandalone_sram5_bus_sel[0]);
	main_genericstandalone_sram5_we[1] <= (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & main_genericstandalone_sram5_bus_we) & main_genericstandalone_sram5_bus_sel[1]);
	main_genericstandalone_sram5_we[2] <= (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & main_genericstandalone_sram5_bus_we) & main_genericstandalone_sram5_bus_sel[2]);
	main_genericstandalone_sram5_we[3] <= (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & main_genericstandalone_sram5_bus_we) & main_genericstandalone_sram5_bus_sel[3]);
	main_genericstandalone_sram5_we[4] <= (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & main_genericstandalone_sram5_bus_we) & main_genericstandalone_sram5_bus_sel[4]);
	main_genericstandalone_sram5_we[5] <= (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & main_genericstandalone_sram5_bus_we) & main_genericstandalone_sram5_bus_sel[5]);
	main_genericstandalone_sram5_we[6] <= (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & main_genericstandalone_sram5_bus_we) & main_genericstandalone_sram5_bus_sel[6]);
	main_genericstandalone_sram5_we[7] <= (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & main_genericstandalone_sram5_bus_we) & main_genericstandalone_sram5_bus_sel[7]);
// synthesis translate_off
	dummy_d_71 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram5_adr = main_genericstandalone_sram5_bus_adr[7:0];
assign main_genericstandalone_sram5_bus_dat_r = main_genericstandalone_sram5_dat_r;
assign main_genericstandalone_sram5_dat_w = main_genericstandalone_sram5_bus_dat_w;

// synthesis translate_off
reg dummy_d_72;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram6_we <= 8'd0;
	main_genericstandalone_sram6_we[0] <= (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & main_genericstandalone_sram6_bus_we) & main_genericstandalone_sram6_bus_sel[0]);
	main_genericstandalone_sram6_we[1] <= (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & main_genericstandalone_sram6_bus_we) & main_genericstandalone_sram6_bus_sel[1]);
	main_genericstandalone_sram6_we[2] <= (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & main_genericstandalone_sram6_bus_we) & main_genericstandalone_sram6_bus_sel[2]);
	main_genericstandalone_sram6_we[3] <= (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & main_genericstandalone_sram6_bus_we) & main_genericstandalone_sram6_bus_sel[3]);
	main_genericstandalone_sram6_we[4] <= (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & main_genericstandalone_sram6_bus_we) & main_genericstandalone_sram6_bus_sel[4]);
	main_genericstandalone_sram6_we[5] <= (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & main_genericstandalone_sram6_bus_we) & main_genericstandalone_sram6_bus_sel[5]);
	main_genericstandalone_sram6_we[6] <= (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & main_genericstandalone_sram6_bus_we) & main_genericstandalone_sram6_bus_sel[6]);
	main_genericstandalone_sram6_we[7] <= (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & main_genericstandalone_sram6_bus_we) & main_genericstandalone_sram6_bus_sel[7]);
// synthesis translate_off
	dummy_d_72 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram6_adr = main_genericstandalone_sram6_bus_adr[7:0];
assign main_genericstandalone_sram6_bus_dat_r = main_genericstandalone_sram6_dat_r;
assign main_genericstandalone_sram6_dat_w = main_genericstandalone_sram6_bus_dat_w;

// synthesis translate_off
reg dummy_d_73;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram7_we <= 8'd0;
	main_genericstandalone_sram7_we[0] <= (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & main_genericstandalone_sram7_bus_we) & main_genericstandalone_sram7_bus_sel[0]);
	main_genericstandalone_sram7_we[1] <= (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & main_genericstandalone_sram7_bus_we) & main_genericstandalone_sram7_bus_sel[1]);
	main_genericstandalone_sram7_we[2] <= (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & main_genericstandalone_sram7_bus_we) & main_genericstandalone_sram7_bus_sel[2]);
	main_genericstandalone_sram7_we[3] <= (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & main_genericstandalone_sram7_bus_we) & main_genericstandalone_sram7_bus_sel[3]);
	main_genericstandalone_sram7_we[4] <= (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & main_genericstandalone_sram7_bus_we) & main_genericstandalone_sram7_bus_sel[4]);
	main_genericstandalone_sram7_we[5] <= (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & main_genericstandalone_sram7_bus_we) & main_genericstandalone_sram7_bus_sel[5]);
	main_genericstandalone_sram7_we[6] <= (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & main_genericstandalone_sram7_bus_we) & main_genericstandalone_sram7_bus_sel[6]);
	main_genericstandalone_sram7_we[7] <= (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & main_genericstandalone_sram7_bus_we) & main_genericstandalone_sram7_bus_sel[7]);
// synthesis translate_off
	dummy_d_73 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram7_adr = main_genericstandalone_sram7_bus_adr[7:0];
assign main_genericstandalone_sram7_bus_dat_r = main_genericstandalone_sram7_dat_r;
assign main_genericstandalone_sram7_dat_w = main_genericstandalone_sram7_bus_dat_w;

// synthesis translate_off
reg dummy_d_74;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_slave_sel <= 8'd0;
	main_genericstandalone_slave_sel[0] <= (main_genericstandalone_bus_bus_adr[10:8] == 1'd0);
	main_genericstandalone_slave_sel[1] <= (main_genericstandalone_bus_bus_adr[10:8] == 1'd1);
	main_genericstandalone_slave_sel[2] <= (main_genericstandalone_bus_bus_adr[10:8] == 2'd2);
	main_genericstandalone_slave_sel[3] <= (main_genericstandalone_bus_bus_adr[10:8] == 2'd3);
	main_genericstandalone_slave_sel[4] <= (main_genericstandalone_bus_bus_adr[10:8] == 3'd4);
	main_genericstandalone_slave_sel[5] <= (main_genericstandalone_bus_bus_adr[10:8] == 3'd5);
	main_genericstandalone_slave_sel[6] <= (main_genericstandalone_bus_bus_adr[10:8] == 3'd6);
	main_genericstandalone_slave_sel[7] <= (main_genericstandalone_bus_bus_adr[10:8] == 3'd7);
// synthesis translate_off
	dummy_d_74 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram0_bus_adr = main_genericstandalone_bus_bus_adr;
assign main_genericstandalone_sram0_bus_dat_w = main_genericstandalone_bus_bus_dat_w;
assign main_genericstandalone_sram0_bus_sel = main_genericstandalone_bus_bus_sel;
assign main_genericstandalone_sram0_bus_stb = main_genericstandalone_bus_bus_stb;
assign main_genericstandalone_sram0_bus_we = main_genericstandalone_bus_bus_we;
assign main_genericstandalone_sram0_bus_cti = main_genericstandalone_bus_bus_cti;
assign main_genericstandalone_sram0_bus_bte = main_genericstandalone_bus_bus_bte;
assign main_genericstandalone_sram1_bus_adr = main_genericstandalone_bus_bus_adr;
assign main_genericstandalone_sram1_bus_dat_w = main_genericstandalone_bus_bus_dat_w;
assign main_genericstandalone_sram1_bus_sel = main_genericstandalone_bus_bus_sel;
assign main_genericstandalone_sram1_bus_stb = main_genericstandalone_bus_bus_stb;
assign main_genericstandalone_sram1_bus_we = main_genericstandalone_bus_bus_we;
assign main_genericstandalone_sram1_bus_cti = main_genericstandalone_bus_bus_cti;
assign main_genericstandalone_sram1_bus_bte = main_genericstandalone_bus_bus_bte;
assign main_genericstandalone_sram2_bus_adr = main_genericstandalone_bus_bus_adr;
assign main_genericstandalone_sram2_bus_dat_w = main_genericstandalone_bus_bus_dat_w;
assign main_genericstandalone_sram2_bus_sel = main_genericstandalone_bus_bus_sel;
assign main_genericstandalone_sram2_bus_stb = main_genericstandalone_bus_bus_stb;
assign main_genericstandalone_sram2_bus_we = main_genericstandalone_bus_bus_we;
assign main_genericstandalone_sram2_bus_cti = main_genericstandalone_bus_bus_cti;
assign main_genericstandalone_sram2_bus_bte = main_genericstandalone_bus_bus_bte;
assign main_genericstandalone_sram3_bus_adr = main_genericstandalone_bus_bus_adr;
assign main_genericstandalone_sram3_bus_dat_w = main_genericstandalone_bus_bus_dat_w;
assign main_genericstandalone_sram3_bus_sel = main_genericstandalone_bus_bus_sel;
assign main_genericstandalone_sram3_bus_stb = main_genericstandalone_bus_bus_stb;
assign main_genericstandalone_sram3_bus_we = main_genericstandalone_bus_bus_we;
assign main_genericstandalone_sram3_bus_cti = main_genericstandalone_bus_bus_cti;
assign main_genericstandalone_sram3_bus_bte = main_genericstandalone_bus_bus_bte;
assign main_genericstandalone_sram4_bus_adr = main_genericstandalone_bus_bus_adr;
assign main_genericstandalone_sram4_bus_dat_w = main_genericstandalone_bus_bus_dat_w;
assign main_genericstandalone_sram4_bus_sel = main_genericstandalone_bus_bus_sel;
assign main_genericstandalone_sram4_bus_stb = main_genericstandalone_bus_bus_stb;
assign main_genericstandalone_sram4_bus_we = main_genericstandalone_bus_bus_we;
assign main_genericstandalone_sram4_bus_cti = main_genericstandalone_bus_bus_cti;
assign main_genericstandalone_sram4_bus_bte = main_genericstandalone_bus_bus_bte;
assign main_genericstandalone_sram5_bus_adr = main_genericstandalone_bus_bus_adr;
assign main_genericstandalone_sram5_bus_dat_w = main_genericstandalone_bus_bus_dat_w;
assign main_genericstandalone_sram5_bus_sel = main_genericstandalone_bus_bus_sel;
assign main_genericstandalone_sram5_bus_stb = main_genericstandalone_bus_bus_stb;
assign main_genericstandalone_sram5_bus_we = main_genericstandalone_bus_bus_we;
assign main_genericstandalone_sram5_bus_cti = main_genericstandalone_bus_bus_cti;
assign main_genericstandalone_sram5_bus_bte = main_genericstandalone_bus_bus_bte;
assign main_genericstandalone_sram6_bus_adr = main_genericstandalone_bus_bus_adr;
assign main_genericstandalone_sram6_bus_dat_w = main_genericstandalone_bus_bus_dat_w;
assign main_genericstandalone_sram6_bus_sel = main_genericstandalone_bus_bus_sel;
assign main_genericstandalone_sram6_bus_stb = main_genericstandalone_bus_bus_stb;
assign main_genericstandalone_sram6_bus_we = main_genericstandalone_bus_bus_we;
assign main_genericstandalone_sram6_bus_cti = main_genericstandalone_bus_bus_cti;
assign main_genericstandalone_sram6_bus_bte = main_genericstandalone_bus_bus_bte;
assign main_genericstandalone_sram7_bus_adr = main_genericstandalone_bus_bus_adr;
assign main_genericstandalone_sram7_bus_dat_w = main_genericstandalone_bus_bus_dat_w;
assign main_genericstandalone_sram7_bus_sel = main_genericstandalone_bus_bus_sel;
assign main_genericstandalone_sram7_bus_stb = main_genericstandalone_bus_bus_stb;
assign main_genericstandalone_sram7_bus_we = main_genericstandalone_bus_bus_we;
assign main_genericstandalone_sram7_bus_cti = main_genericstandalone_bus_bus_cti;
assign main_genericstandalone_sram7_bus_bte = main_genericstandalone_bus_bus_bte;
assign main_genericstandalone_sram0_bus_cyc = (main_genericstandalone_bus_bus_cyc & main_genericstandalone_slave_sel[0]);
assign main_genericstandalone_sram1_bus_cyc = (main_genericstandalone_bus_bus_cyc & main_genericstandalone_slave_sel[1]);
assign main_genericstandalone_sram2_bus_cyc = (main_genericstandalone_bus_bus_cyc & main_genericstandalone_slave_sel[2]);
assign main_genericstandalone_sram3_bus_cyc = (main_genericstandalone_bus_bus_cyc & main_genericstandalone_slave_sel[3]);
assign main_genericstandalone_sram4_bus_cyc = (main_genericstandalone_bus_bus_cyc & main_genericstandalone_slave_sel[4]);
assign main_genericstandalone_sram5_bus_cyc = (main_genericstandalone_bus_bus_cyc & main_genericstandalone_slave_sel[5]);
assign main_genericstandalone_sram6_bus_cyc = (main_genericstandalone_bus_bus_cyc & main_genericstandalone_slave_sel[6]);
assign main_genericstandalone_sram7_bus_cyc = (main_genericstandalone_bus_bus_cyc & main_genericstandalone_slave_sel[7]);
assign main_genericstandalone_bus_bus_ack = (((((((main_genericstandalone_sram0_bus_ack | main_genericstandalone_sram1_bus_ack) | main_genericstandalone_sram2_bus_ack) | main_genericstandalone_sram3_bus_ack) | main_genericstandalone_sram4_bus_ack) | main_genericstandalone_sram5_bus_ack) | main_genericstandalone_sram6_bus_ack) | main_genericstandalone_sram7_bus_ack);
assign main_genericstandalone_bus_bus_err = (((((((main_genericstandalone_sram0_bus_err | main_genericstandalone_sram1_bus_err) | main_genericstandalone_sram2_bus_err) | main_genericstandalone_sram3_bus_err) | main_genericstandalone_sram4_bus_err) | main_genericstandalone_sram5_bus_err) | main_genericstandalone_sram6_bus_err) | main_genericstandalone_sram7_bus_err);
assign main_genericstandalone_bus_bus_dat_r = (((((((({64{main_genericstandalone_slave_sel_r[0]}} & main_genericstandalone_sram0_bus_dat_r) | ({64{main_genericstandalone_slave_sel_r[1]}} & main_genericstandalone_sram1_bus_dat_r)) | ({64{main_genericstandalone_slave_sel_r[2]}} & main_genericstandalone_sram2_bus_dat_r)) | ({64{main_genericstandalone_slave_sel_r[3]}} & main_genericstandalone_sram3_bus_dat_r)) | ({64{main_genericstandalone_slave_sel_r[4]}} & main_genericstandalone_sram4_bus_dat_r)) | ({64{main_genericstandalone_slave_sel_r[5]}} & main_genericstandalone_sram5_bus_dat_r)) | ({64{main_genericstandalone_slave_sel_r[6]}} & main_genericstandalone_sram6_bus_dat_r)) | ({64{main_genericstandalone_slave_sel_r[7]}} & main_genericstandalone_sram7_bus_dat_r));
assign sys_kernel_clk = sys_clk;
assign sys_kernel_rst = main_genericstandalone_kernel_cpu_storage;
assign builder_shared_adr = builder_comb_rhs_self0;
assign builder_shared_dat_w = builder_comb_rhs_self1;
assign builder_shared_sel = builder_comb_rhs_self2;
assign builder_shared_cyc = builder_comb_rhs_self3;
assign builder_shared_stb = builder_comb_rhs_self4;
assign builder_shared_we = builder_comb_rhs_self5;
assign builder_shared_cti = builder_comb_rhs_self6;
assign builder_shared_bte = builder_comb_rhs_self7;
assign main_genericstandalone_kernel_cpu_ibus_dat_r = builder_shared_dat_r;
assign main_genericstandalone_kernel_cpu_dbus_dat_r = builder_shared_dat_r;
assign main_genericstandalone_kernel_cpu_ibus_ack = (builder_shared_ack & (builder_grant == 1'd0));
assign main_genericstandalone_kernel_cpu_dbus_ack = (builder_shared_ack & (builder_grant == 1'd1));
assign main_genericstandalone_kernel_cpu_ibus_err = (builder_shared_err & (builder_grant == 1'd0));
assign main_genericstandalone_kernel_cpu_dbus_err = (builder_shared_err & (builder_grant == 1'd1));
assign builder_request = {(main_genericstandalone_kernel_cpu_dbus_cyc & (~(main_genericstandalone_kernel_cpu_dbus_ack & (main_genericstandalone_kernel_cpu_dbus_cti != 2'd2)))), (main_genericstandalone_kernel_cpu_ibus_cyc & (~(main_genericstandalone_kernel_cpu_ibus_ack & (main_genericstandalone_kernel_cpu_ibus_cti != 2'd2))))};

// synthesis translate_off
reg dummy_d_75;
// synthesis translate_on
always @(*) begin
	builder_slave_sel <= 5'd0;
	builder_slave_sel[0] <= ((1'd1 & (~builder_shared_adr[26])) & builder_shared_adr[27]);
	builder_slave_sel[1] <= ((1'd1 & builder_shared_adr[26]) & builder_shared_adr[27]);
	builder_slave_sel[2] <= (((1'd1 & (~builder_shared_adr[25])) & (~builder_shared_adr[27])) & builder_shared_adr[26]);
	builder_slave_sel[3] <= (((1'd1 & (~builder_shared_adr[27])) & builder_shared_adr[25]) & builder_shared_adr[26]);
	builder_slave_sel[4] <= ((1'd1 & (~builder_shared_adr[26])) & (~builder_shared_adr[27]));
// synthesis translate_off
	dummy_d_75 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_kernel_cpu_wb_sdram_adr = builder_shared_adr;
assign main_genericstandalone_kernel_cpu_wb_sdram_dat_w = builder_shared_dat_w;
assign main_genericstandalone_kernel_cpu_wb_sdram_sel = builder_shared_sel;
assign main_genericstandalone_kernel_cpu_wb_sdram_stb = builder_shared_stb;
assign main_genericstandalone_kernel_cpu_wb_sdram_we = builder_shared_we;
assign main_genericstandalone_kernel_cpu_wb_sdram_cti = builder_shared_cti;
assign main_genericstandalone_kernel_cpu_wb_sdram_bte = builder_shared_bte;
assign main_genericstandalone_mailbox_i2_adr = builder_shared_adr;
assign main_genericstandalone_mailbox_i2_dat_w = builder_shared_dat_w;
assign main_genericstandalone_mailbox_i2_sel = builder_shared_sel;
assign main_genericstandalone_mailbox_i2_stb = builder_shared_stb;
assign main_genericstandalone_mailbox_i2_we = builder_shared_we;
assign main_genericstandalone_mailbox_i2_cti = builder_shared_cti;
assign main_genericstandalone_mailbox_i2_bte = builder_shared_bte;
assign main_genericstandalone_interface0_csr_bus_adr = builder_shared_adr;
assign main_genericstandalone_interface0_csr_bus_dat_w = builder_shared_dat_w;
assign main_genericstandalone_interface0_csr_bus_sel = builder_shared_sel;
assign main_genericstandalone_interface0_csr_bus_stb = builder_shared_stb;
assign main_genericstandalone_interface0_csr_bus_we = builder_shared_we;
assign main_genericstandalone_interface0_csr_bus_cti = builder_shared_cti;
assign main_genericstandalone_interface0_csr_bus_bte = builder_shared_bte;
assign main_genericstandalone_interface1_csr_bus_adr = builder_shared_adr;
assign main_genericstandalone_interface1_csr_bus_dat_w = builder_shared_dat_w;
assign main_genericstandalone_interface1_csr_bus_sel = builder_shared_sel;
assign main_genericstandalone_interface1_csr_bus_stb = builder_shared_stb;
assign main_genericstandalone_interface1_csr_bus_we = builder_shared_we;
assign main_genericstandalone_interface1_csr_bus_cti = builder_shared_cti;
assign main_genericstandalone_interface1_csr_bus_bte = builder_shared_bte;
assign main_genericstandalone_interface2_csr_bus_adr = builder_shared_adr;
assign main_genericstandalone_interface2_csr_bus_dat_w = builder_shared_dat_w;
assign main_genericstandalone_interface2_csr_bus_sel = builder_shared_sel;
assign main_genericstandalone_interface2_csr_bus_stb = builder_shared_stb;
assign main_genericstandalone_interface2_csr_bus_we = builder_shared_we;
assign main_genericstandalone_interface2_csr_bus_cti = builder_shared_cti;
assign main_genericstandalone_interface2_csr_bus_bte = builder_shared_bte;
assign main_genericstandalone_kernel_cpu_wb_sdram_cyc = (builder_shared_cyc & builder_slave_sel[0]);
assign main_genericstandalone_mailbox_i2_cyc = (builder_shared_cyc & builder_slave_sel[1]);
assign main_genericstandalone_interface0_csr_bus_cyc = (builder_shared_cyc & builder_slave_sel[2]);
assign main_genericstandalone_interface1_csr_bus_cyc = (builder_shared_cyc & builder_slave_sel[3]);
assign main_genericstandalone_interface2_csr_bus_cyc = (builder_shared_cyc & builder_slave_sel[4]);
assign builder_shared_ack = ((((main_genericstandalone_kernel_cpu_wb_sdram_ack | main_genericstandalone_mailbox_i2_ack) | main_genericstandalone_interface0_csr_bus_ack) | main_genericstandalone_interface1_csr_bus_ack) | main_genericstandalone_interface2_csr_bus_ack);
assign builder_shared_err = ((((main_genericstandalone_kernel_cpu_wb_sdram_err | main_genericstandalone_mailbox_i2_err) | main_genericstandalone_interface0_csr_bus_err) | main_genericstandalone_interface1_csr_bus_err) | main_genericstandalone_interface2_csr_bus_err);
assign builder_shared_dat_r = ((((({64{builder_slave_sel_r[0]}} & main_genericstandalone_kernel_cpu_wb_sdram_dat_r) | ({64{builder_slave_sel_r[1]}} & main_genericstandalone_mailbox_i2_dat_r)) | ({64{builder_slave_sel_r[2]}} & main_genericstandalone_interface0_csr_bus_dat_r)) | ({64{builder_slave_sel_r[3]}} & main_genericstandalone_interface1_csr_bus_dat_r)) | ({64{builder_slave_sel_r[4]}} & main_genericstandalone_interface2_csr_bus_dat_r));
assign {error_led} = main_genericstandalone_error_led_storage;
assign main_genericstandalone_i2c_tstriple0_o = main_genericstandalone_i2c_out_storage[0];
assign main_genericstandalone_i2c_tstriple0_oe = main_genericstandalone_i2c_oe_storage[0];

// synthesis translate_off
reg dummy_d_76;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_i2c_status0 <= 2'd0;
	main_genericstandalone_i2c_status0[0] <= main_genericstandalone_i2c_status1;
	main_genericstandalone_i2c_status0[1] <= main_genericstandalone_i2c_status2;
// synthesis translate_off
	dummy_d_76 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_i2c_tstriple1_o = main_genericstandalone_i2c_out_storage[1];
assign main_genericstandalone_i2c_tstriple1_oe = main_genericstandalone_i2c_oe_storage[1];
assign main_inout_8x0_serdes_oe = main_inout_8x0_inout_8x0_oe;
assign main_inout_8x0_inout_8x0_input_state = main_inout_8x0_serdes_i0[7];
assign main_inout_8x0_inout_8x0_i = ((main_inout_8x0_serdes_i0 ^ {main_inout_8x0_serdes_i0, main_inout_8x0_inout_8x0_i_d}) & ((main_inout_8x0_serdes_i0 & {8{main_inout_8x0_inout_8x0_sensitivity[0]}}) | ((~main_inout_8x0_serdes_i0) & {8{main_inout_8x0_inout_8x0_sensitivity[1]}})));
assign main_inout_8x0_serdes_i0 = main_inout_8x0_serdes_i1;
assign main_inout_8x0_serdes_o1 = main_inout_8x0_serdes_o0;
assign main_inout_8x0_serdes_t_in = (~main_inout_8x0_serdes_oe);

// synthesis translate_off
reg dummy_d_77;
// synthesis translate_on
always @(*) begin
	main_inout_8x0_inout_8x0_o <= 3'd0;
	if (main_inout_8x0_inout_8x0_i[7]) begin
		main_inout_8x0_inout_8x0_o <= 3'd7;
	end
	if (main_inout_8x0_inout_8x0_i[6]) begin
		main_inout_8x0_inout_8x0_o <= 3'd6;
	end
	if (main_inout_8x0_inout_8x0_i[5]) begin
		main_inout_8x0_inout_8x0_o <= 3'd5;
	end
	if (main_inout_8x0_inout_8x0_i[4]) begin
		main_inout_8x0_inout_8x0_o <= 3'd4;
	end
	if (main_inout_8x0_inout_8x0_i[3]) begin
		main_inout_8x0_inout_8x0_o <= 2'd3;
	end
	if (main_inout_8x0_inout_8x0_i[2]) begin
		main_inout_8x0_inout_8x0_o <= 2'd2;
	end
	if (main_inout_8x0_inout_8x0_i[1]) begin
		main_inout_8x0_inout_8x0_o <= 1'd1;
	end
	if (main_inout_8x0_inout_8x0_i[0]) begin
		main_inout_8x0_inout_8x0_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_77 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x0_inout_8x0_n = (main_inout_8x0_inout_8x0_i == 1'd0);
assign main_inout_8x1_serdes_oe = main_inout_8x1_inout_8x1_oe;
assign main_inout_8x1_inout_8x1_input_state = main_inout_8x1_serdes_i0[7];
assign main_inout_8x1_inout_8x1_i = ((main_inout_8x1_serdes_i0 ^ {main_inout_8x1_serdes_i0, main_inout_8x1_inout_8x1_i_d}) & ((main_inout_8x1_serdes_i0 & {8{main_inout_8x1_inout_8x1_sensitivity[0]}}) | ((~main_inout_8x1_serdes_i0) & {8{main_inout_8x1_inout_8x1_sensitivity[1]}})));
assign main_inout_8x1_serdes_i0 = main_inout_8x1_serdes_i1;
assign main_inout_8x1_serdes_o1 = main_inout_8x1_serdes_o0;
assign main_inout_8x1_serdes_t_in = (~main_inout_8x1_serdes_oe);

// synthesis translate_off
reg dummy_d_78;
// synthesis translate_on
always @(*) begin
	main_inout_8x1_inout_8x1_o <= 3'd0;
	if (main_inout_8x1_inout_8x1_i[7]) begin
		main_inout_8x1_inout_8x1_o <= 3'd7;
	end
	if (main_inout_8x1_inout_8x1_i[6]) begin
		main_inout_8x1_inout_8x1_o <= 3'd6;
	end
	if (main_inout_8x1_inout_8x1_i[5]) begin
		main_inout_8x1_inout_8x1_o <= 3'd5;
	end
	if (main_inout_8x1_inout_8x1_i[4]) begin
		main_inout_8x1_inout_8x1_o <= 3'd4;
	end
	if (main_inout_8x1_inout_8x1_i[3]) begin
		main_inout_8x1_inout_8x1_o <= 2'd3;
	end
	if (main_inout_8x1_inout_8x1_i[2]) begin
		main_inout_8x1_inout_8x1_o <= 2'd2;
	end
	if (main_inout_8x1_inout_8x1_i[1]) begin
		main_inout_8x1_inout_8x1_o <= 1'd1;
	end
	if (main_inout_8x1_inout_8x1_i[0]) begin
		main_inout_8x1_inout_8x1_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_78 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x1_inout_8x1_n = (main_inout_8x1_inout_8x1_i == 1'd0);
assign main_inout_8x2_serdes_oe = main_inout_8x2_inout_8x2_oe;
assign main_inout_8x2_inout_8x2_input_state = main_inout_8x2_serdes_i0[7];
assign main_inout_8x2_inout_8x2_i = ((main_inout_8x2_serdes_i0 ^ {main_inout_8x2_serdes_i0, main_inout_8x2_inout_8x2_i_d}) & ((main_inout_8x2_serdes_i0 & {8{main_inout_8x2_inout_8x2_sensitivity[0]}}) | ((~main_inout_8x2_serdes_i0) & {8{main_inout_8x2_inout_8x2_sensitivity[1]}})));
assign main_inout_8x2_serdes_i0 = main_inout_8x2_serdes_i1;
assign main_inout_8x2_serdes_o1 = main_inout_8x2_serdes_o0;
assign main_inout_8x2_serdes_t_in = (~main_inout_8x2_serdes_oe);

// synthesis translate_off
reg dummy_d_79;
// synthesis translate_on
always @(*) begin
	main_inout_8x2_inout_8x2_o <= 3'd0;
	if (main_inout_8x2_inout_8x2_i[7]) begin
		main_inout_8x2_inout_8x2_o <= 3'd7;
	end
	if (main_inout_8x2_inout_8x2_i[6]) begin
		main_inout_8x2_inout_8x2_o <= 3'd6;
	end
	if (main_inout_8x2_inout_8x2_i[5]) begin
		main_inout_8x2_inout_8x2_o <= 3'd5;
	end
	if (main_inout_8x2_inout_8x2_i[4]) begin
		main_inout_8x2_inout_8x2_o <= 3'd4;
	end
	if (main_inout_8x2_inout_8x2_i[3]) begin
		main_inout_8x2_inout_8x2_o <= 2'd3;
	end
	if (main_inout_8x2_inout_8x2_i[2]) begin
		main_inout_8x2_inout_8x2_o <= 2'd2;
	end
	if (main_inout_8x2_inout_8x2_i[1]) begin
		main_inout_8x2_inout_8x2_o <= 1'd1;
	end
	if (main_inout_8x2_inout_8x2_i[0]) begin
		main_inout_8x2_inout_8x2_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_79 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x2_inout_8x2_n = (main_inout_8x2_inout_8x2_i == 1'd0);
assign main_inout_8x3_serdes_oe = main_inout_8x3_inout_8x3_oe;
assign main_inout_8x3_inout_8x3_input_state = main_inout_8x3_serdes_i0[7];
assign main_inout_8x3_inout_8x3_i = ((main_inout_8x3_serdes_i0 ^ {main_inout_8x3_serdes_i0, main_inout_8x3_inout_8x3_i_d}) & ((main_inout_8x3_serdes_i0 & {8{main_inout_8x3_inout_8x3_sensitivity[0]}}) | ((~main_inout_8x3_serdes_i0) & {8{main_inout_8x3_inout_8x3_sensitivity[1]}})));
assign main_inout_8x3_serdes_i0 = main_inout_8x3_serdes_i1;
assign main_inout_8x3_serdes_o1 = main_inout_8x3_serdes_o0;
assign main_inout_8x3_serdes_t_in = (~main_inout_8x3_serdes_oe);

// synthesis translate_off
reg dummy_d_80;
// synthesis translate_on
always @(*) begin
	main_inout_8x3_inout_8x3_o <= 3'd0;
	if (main_inout_8x3_inout_8x3_i[7]) begin
		main_inout_8x3_inout_8x3_o <= 3'd7;
	end
	if (main_inout_8x3_inout_8x3_i[6]) begin
		main_inout_8x3_inout_8x3_o <= 3'd6;
	end
	if (main_inout_8x3_inout_8x3_i[5]) begin
		main_inout_8x3_inout_8x3_o <= 3'd5;
	end
	if (main_inout_8x3_inout_8x3_i[4]) begin
		main_inout_8x3_inout_8x3_o <= 3'd4;
	end
	if (main_inout_8x3_inout_8x3_i[3]) begin
		main_inout_8x3_inout_8x3_o <= 2'd3;
	end
	if (main_inout_8x3_inout_8x3_i[2]) begin
		main_inout_8x3_inout_8x3_o <= 2'd2;
	end
	if (main_inout_8x3_inout_8x3_i[1]) begin
		main_inout_8x3_inout_8x3_o <= 1'd1;
	end
	if (main_inout_8x3_inout_8x3_i[0]) begin
		main_inout_8x3_inout_8x3_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_80 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x3_inout_8x3_n = (main_inout_8x3_inout_8x3_i == 1'd0);
assign main_spimaster0_spimachine0_length0 = main_spimaster0_config_length0;
assign main_spimaster0_spimachine0_end0 = main_spimaster0_config_end0;
assign main_spimaster0_spimachine0_div0 = main_spimaster0_config_div0;
assign main_spimaster0_spimachine0_clk_phase0 = main_spimaster0_config_clk_phase0;
assign main_spimaster0_spimachine0_lsb_first0 = main_spimaster0_config_lsb_first0;
assign main_spimaster0_interface_half_duplex0 = main_spimaster0_config_half_duplex0;
assign main_spimaster0_interface_cs0 = main_spimaster0_config_cs0;
assign main_spimaster0_interface_cs_polarity0 = {3{main_spimaster0_config_cs_polarity0}};
assign main_spimaster0_interface_clk_polarity0 = main_spimaster0_config_clk_polarity0;
assign main_spimaster0_interface_offline0 = main_spimaster0_config_offline0;
assign main_spimaster0_interface_cs_next0 = main_spimaster0_spimachine0_cs_next0;
assign main_spimaster0_interface_clk_next0 = main_spimaster0_spimachine0_clk_next0;
assign main_spimaster0_interface_ce0 = main_spimaster0_spimachine0_ce0;
assign main_spimaster0_interface_sample0 = main_spimaster0_spimachine0_sample0;
assign main_spimaster0_spimachine0_sdi0 = main_spimaster0_interface_sdi0;
assign main_spimaster0_interface_sdo0 = main_spimaster0_spimachine0_sdo0;
assign main_spimaster0_spimachine0_load0 = ((main_spimaster0_ointerface0_stb0 & main_spimaster0_spimachine0_writable0) & (~main_spimaster0_ointerface0_address0));
assign main_spimaster0_spimachine0_pdo0 = main_spimaster0_ointerface0_data0;
assign main_spimaster0_ointerface0_busy0 = (~main_spimaster0_spimachine0_writable0);
assign main_spimaster0_iinterface0_stb0 = (main_spimaster0_spimachine0_readable0 & main_spimaster0_read0);
assign main_spimaster0_iinterface0_data0 = main_spimaster0_spimachine0_pdi0;
assign main_spimaster0_interface_sdi0 = (main_spimaster0_interface_half_duplex0 ? main_spimaster0_interface_mosi_reg0 : main_spimaster0_interface_miso_reg0);
assign main_spimaster0_spimachine0_ce0 = (main_spimaster0_spimachine0_done0 & main_spimaster0_spimachine0_count0);
assign main_spimaster0_spimachine0_pdi0 = (main_spimaster0_spimachine0_lsb_first0 ? {main_spimaster0_spimachine0_sdi0, main_spimaster0_spimachine0_sr0[31:1]} : {main_spimaster0_spimachine0_sr0[30:0], main_spimaster0_spimachine0_sdi0});
assign main_spimaster0_spimachine0_cnt_done0 = (main_spimaster0_spimachine0_cnt0 == 1'd0);
assign main_spimaster0_spimachine0_done0 = (main_spimaster0_spimachine0_cnt_done0 & (~main_spimaster0_spimachine0_do_extend0));

// synthesis translate_off
reg dummy_d_81;
// synthesis translate_on
always @(*) begin
	main_spimaster0_spimachine0_clk_next0 <= 1'd0;
	main_spimaster0_spimachine0_cs_next0 <= 1'd0;
	main_spimaster0_spimachine0_idle0 <= 1'd0;
	main_spimaster0_spimachine0_readable0 <= 1'd0;
	main_spimaster0_spimachine0_writable0 <= 1'd0;
	main_spimaster0_spimachine0_load1 <= 1'd0;
	main_spimaster0_spimachine0_shift0 <= 1'd0;
	main_spimaster0_spimachine0_sample0 <= 1'd0;
	main_spimaster0_spimachine0_extend0 <= 1'd0;
	main_spimaster0_spimachine0_count0 <= 1'd0;
	builder_spimaster0_next_state <= 3'd0;
	builder_spimaster0_next_state <= builder_spimaster0_state;
	case (builder_spimaster0_state)
		1'd1: begin
			main_spimaster0_spimachine0_cs_next0 <= 1'd1;
			main_spimaster0_spimachine0_count0 <= 1'd1;
			main_spimaster0_spimachine0_extend0 <= 1'd1;
			main_spimaster0_spimachine0_clk_next0 <= 1'd1;
			if (main_spimaster0_spimachine0_done0) begin
				builder_spimaster0_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster0_spimachine0_cs_next0 <= 1'd1;
			main_spimaster0_spimachine0_count0 <= 1'd1;
			main_spimaster0_spimachine0_clk_next0 <= (~main_spimaster0_spimachine0_clk_phase0);
			if (main_spimaster0_spimachine0_done0) begin
				main_spimaster0_spimachine0_sample0 <= 1'd1;
				builder_spimaster0_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster0_spimachine0_cs_next0 <= 1'd1;
			main_spimaster0_spimachine0_count0 <= 1'd1;
			main_spimaster0_spimachine0_extend0 <= 1'd1;
			main_spimaster0_spimachine0_clk_next0 <= main_spimaster0_spimachine0_clk_phase0;
			if (main_spimaster0_spimachine0_done0) begin
				if ((main_spimaster0_spimachine0_n0 == 1'd0)) begin
					main_spimaster0_spimachine0_readable0 <= 1'd1;
					main_spimaster0_spimachine0_writable0 <= 1'd1;
					if (main_spimaster0_spimachine0_end1) begin
						main_spimaster0_spimachine0_clk_next0 <= 1'd0;
						main_spimaster0_spimachine0_writable0 <= 1'd0;
						if (main_spimaster0_spimachine0_clk_phase0) begin
							main_spimaster0_spimachine0_cs_next0 <= 1'd0;
							builder_spimaster0_next_state <= 3'd5;
						end else begin
							builder_spimaster0_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster0_spimachine0_load0) begin
							main_spimaster0_spimachine0_load1 <= 1'd1;
							builder_spimaster0_next_state <= 2'd2;
						end else begin
							main_spimaster0_spimachine0_count0 <= 1'd0;
						end
					end
				end else begin
					main_spimaster0_spimachine0_shift0 <= 1'd1;
					builder_spimaster0_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster0_spimachine0_count0 <= 1'd1;
			if (main_spimaster0_spimachine0_done0) begin
				builder_spimaster0_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster0_spimachine0_done0) begin
				builder_spimaster0_next_state <= 1'd0;
			end else begin
				main_spimaster0_spimachine0_count0 <= 1'd1;
			end
		end
		default: begin
			main_spimaster0_spimachine0_idle0 <= 1'd1;
			main_spimaster0_spimachine0_writable0 <= 1'd1;
			main_spimaster0_spimachine0_cs_next0 <= 1'd1;
			if (main_spimaster0_spimachine0_load0) begin
				main_spimaster0_spimachine0_count0 <= 1'd1;
				main_spimaster0_spimachine0_load1 <= 1'd1;
				if (main_spimaster0_spimachine0_clk_phase0) begin
					builder_spimaster0_next_state <= 1'd1;
				end else begin
					main_spimaster0_spimachine0_extend0 <= 1'd1;
					builder_spimaster0_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_81 <= dummy_s;
// synthesis translate_on
end
assign main_urukulmonitor0_ch_sel0 = (((main_urukulmonitor0_cs == 2'd3) | (main_urukulmonitor0_cs == 3'd4)) & (main_urukulmonitor0_current_address == 1'd0));
assign main_urukulmonitor0_ch_sel1 = (((main_urukulmonitor0_cs == 2'd3) | (main_urukulmonitor0_cs == 3'd5)) & (main_urukulmonitor0_current_address == 1'd0));
assign main_urukulmonitor0_ch_sel2 = (((main_urukulmonitor0_cs == 2'd3) | (main_urukulmonitor0_cs == 3'd6)) & (main_urukulmonitor0_current_address == 1'd0));
assign main_urukulmonitor0_ch_sel3 = (((main_urukulmonitor0_cs == 2'd3) | (main_urukulmonitor0_cs == 3'd7)) & (main_urukulmonitor0_current_address == 1'd0));

// synthesis translate_off
reg dummy_d_82;
// synthesis translate_on
always @(*) begin
	builder_ad9910monitor0_next_state <= 1'd0;
	builder_ad9910monitor0_next_value <= 16'd0;
	builder_ad9910monitor0_next_value_ce <= 1'd0;
	main_urukulmonitor0_ftw0_ad9910monitor0_next_value <= 32'd0;
	main_urukulmonitor0_ftw0_ad9910monitor0_next_value_ce <= 1'd0;
	builder_ad9910monitor0_next_state <= builder_ad9910monitor0_state;
	case (builder_ad9910monitor0_state)
		1'd1: begin
			if (main_urukulmonitor0_ch_sel0) begin
				if ((main_urukulmonitor0_flags & 2'd2)) begin
					main_urukulmonitor0_ftw0_ad9910monitor0_next_value <= main_urukulmonitor0_current_data;
					main_urukulmonitor0_ftw0_ad9910monitor0_next_value_ce <= 1'd1;
					builder_ad9910monitor0_next_state <= 1'd0;
				end
			end
		end
		default: begin
			if ((main_urukulmonitor0_ch_sel0 & (~main_urukulmonitor0_current_data[31]))) begin
				if ((((main_urukulmonitor0_data_length == 4'd8) & (main_urukulmonitor0_current_data[28:24] <= 5'd21)) & (main_urukulmonitor0_current_data[28:24] >= 4'd14))) begin
					builder_ad9910monitor0_next_state <= 1'd1;
				end else begin
					if ((main_urukulmonitor0_current_data[28:24] == 3'd7)) begin
						if (((main_urukulmonitor0_data_length == 5'd24) & (main_urukulmonitor0_flags & 2'd2))) begin
							builder_ad9910monitor0_next_value <= main_urukulmonitor0_current_data[23:8];
							builder_ad9910monitor0_next_value_ce <= 1'd1;
						end else begin
							if ((main_urukulmonitor0_data_length == 4'd8)) begin
								builder_ad9910monitor0_next_state <= 1'd1;
							end
						end
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_82 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_83;
// synthesis translate_on
always @(*) begin
	builder_ad9910monitor1_next_state <= 1'd0;
	builder_ad9910monitor1_next_value <= 16'd0;
	builder_ad9910monitor1_next_value_ce <= 1'd0;
	main_urukulmonitor0_ftw1_ad9910monitor1_next_value <= 32'd0;
	main_urukulmonitor0_ftw1_ad9910monitor1_next_value_ce <= 1'd0;
	builder_ad9910monitor1_next_state <= builder_ad9910monitor1_state;
	case (builder_ad9910monitor1_state)
		1'd1: begin
			if (main_urukulmonitor0_ch_sel1) begin
				if ((main_urukulmonitor0_flags & 2'd2)) begin
					main_urukulmonitor0_ftw1_ad9910monitor1_next_value <= main_urukulmonitor0_current_data;
					main_urukulmonitor0_ftw1_ad9910monitor1_next_value_ce <= 1'd1;
					builder_ad9910monitor1_next_state <= 1'd0;
				end
			end
		end
		default: begin
			if ((main_urukulmonitor0_ch_sel1 & (~main_urukulmonitor0_current_data[31]))) begin
				if ((((main_urukulmonitor0_data_length == 4'd8) & (main_urukulmonitor0_current_data[28:24] <= 5'd21)) & (main_urukulmonitor0_current_data[28:24] >= 4'd14))) begin
					builder_ad9910monitor1_next_state <= 1'd1;
				end else begin
					if ((main_urukulmonitor0_current_data[28:24] == 3'd7)) begin
						if (((main_urukulmonitor0_data_length == 5'd24) & (main_urukulmonitor0_flags & 2'd2))) begin
							builder_ad9910monitor1_next_value <= main_urukulmonitor0_current_data[23:8];
							builder_ad9910monitor1_next_value_ce <= 1'd1;
						end else begin
							if ((main_urukulmonitor0_data_length == 4'd8)) begin
								builder_ad9910monitor1_next_state <= 1'd1;
							end
						end
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_83 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_84;
// synthesis translate_on
always @(*) begin
	builder_ad9910monitor2_next_state <= 1'd0;
	builder_ad9910monitor2_next_value <= 16'd0;
	builder_ad9910monitor2_next_value_ce <= 1'd0;
	main_urukulmonitor0_ftw2_ad9910monitor2_next_value <= 32'd0;
	main_urukulmonitor0_ftw2_ad9910monitor2_next_value_ce <= 1'd0;
	builder_ad9910monitor2_next_state <= builder_ad9910monitor2_state;
	case (builder_ad9910monitor2_state)
		1'd1: begin
			if (main_urukulmonitor0_ch_sel2) begin
				if ((main_urukulmonitor0_flags & 2'd2)) begin
					main_urukulmonitor0_ftw2_ad9910monitor2_next_value <= main_urukulmonitor0_current_data;
					main_urukulmonitor0_ftw2_ad9910monitor2_next_value_ce <= 1'd1;
					builder_ad9910monitor2_next_state <= 1'd0;
				end
			end
		end
		default: begin
			if ((main_urukulmonitor0_ch_sel2 & (~main_urukulmonitor0_current_data[31]))) begin
				if ((((main_urukulmonitor0_data_length == 4'd8) & (main_urukulmonitor0_current_data[28:24] <= 5'd21)) & (main_urukulmonitor0_current_data[28:24] >= 4'd14))) begin
					builder_ad9910monitor2_next_state <= 1'd1;
				end else begin
					if ((main_urukulmonitor0_current_data[28:24] == 3'd7)) begin
						if (((main_urukulmonitor0_data_length == 5'd24) & (main_urukulmonitor0_flags & 2'd2))) begin
							builder_ad9910monitor2_next_value <= main_urukulmonitor0_current_data[23:8];
							builder_ad9910monitor2_next_value_ce <= 1'd1;
						end else begin
							if ((main_urukulmonitor0_data_length == 4'd8)) begin
								builder_ad9910monitor2_next_state <= 1'd1;
							end
						end
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_84 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_85;
// synthesis translate_on
always @(*) begin
	builder_ad9910monitor3_next_state <= 1'd0;
	builder_ad9910monitor3_next_value <= 16'd0;
	builder_ad9910monitor3_next_value_ce <= 1'd0;
	main_urukulmonitor0_ftw3_ad9910monitor3_next_value <= 32'd0;
	main_urukulmonitor0_ftw3_ad9910monitor3_next_value_ce <= 1'd0;
	builder_ad9910monitor3_next_state <= builder_ad9910monitor3_state;
	case (builder_ad9910monitor3_state)
		1'd1: begin
			if (main_urukulmonitor0_ch_sel3) begin
				if ((main_urukulmonitor0_flags & 2'd2)) begin
					main_urukulmonitor0_ftw3_ad9910monitor3_next_value <= main_urukulmonitor0_current_data;
					main_urukulmonitor0_ftw3_ad9910monitor3_next_value_ce <= 1'd1;
					builder_ad9910monitor3_next_state <= 1'd0;
				end
			end
		end
		default: begin
			if ((main_urukulmonitor0_ch_sel3 & (~main_urukulmonitor0_current_data[31]))) begin
				if ((((main_urukulmonitor0_data_length == 4'd8) & (main_urukulmonitor0_current_data[28:24] <= 5'd21)) & (main_urukulmonitor0_current_data[28:24] >= 4'd14))) begin
					builder_ad9910monitor3_next_state <= 1'd1;
				end else begin
					if ((main_urukulmonitor0_current_data[28:24] == 3'd7)) begin
						if (((main_urukulmonitor0_data_length == 5'd24) & (main_urukulmonitor0_flags & 2'd2))) begin
							builder_ad9910monitor3_next_value <= main_urukulmonitor0_current_data[23:8];
							builder_ad9910monitor3_next_value_ce <= 1'd1;
						end else begin
							if ((main_urukulmonitor0_data_length == 4'd8)) begin
								builder_ad9910monitor3_next_state <= 1'd1;
							end
						end
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_85 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster1_spimachine1_length0 = main_spimaster1_config_length0;
assign main_spimaster1_spimachine1_end0 = main_spimaster1_config_end0;
assign main_spimaster1_spimachine1_div0 = main_spimaster1_config_div0;
assign main_spimaster1_spimachine1_clk_phase0 = main_spimaster1_config_clk_phase0;
assign main_spimaster1_spimachine1_lsb_first0 = main_spimaster1_config_lsb_first0;
assign main_spimaster1_interface_half_duplex0 = main_spimaster1_config_half_duplex0;
assign main_spimaster1_interface_cs0 = main_spimaster1_config_cs0;
assign main_spimaster1_interface_cs_polarity0 = {3{main_spimaster1_config_cs_polarity0}};
assign main_spimaster1_interface_clk_polarity0 = main_spimaster1_config_clk_polarity0;
assign main_spimaster1_interface_offline0 = main_spimaster1_config_offline0;
assign main_spimaster1_interface_cs_next0 = main_spimaster1_spimachine1_cs_next0;
assign main_spimaster1_interface_clk_next0 = main_spimaster1_spimachine1_clk_next0;
assign main_spimaster1_interface_ce0 = main_spimaster1_spimachine1_ce0;
assign main_spimaster1_interface_sample0 = main_spimaster1_spimachine1_sample0;
assign main_spimaster1_spimachine1_sdi0 = main_spimaster1_interface_sdi0;
assign main_spimaster1_interface_sdo0 = main_spimaster1_spimachine1_sdo0;
assign main_spimaster1_spimachine1_load0 = ((main_spimaster1_ointerface1_stb0 & main_spimaster1_spimachine1_writable0) & (~main_spimaster1_ointerface1_address0));
assign main_spimaster1_spimachine1_pdo0 = main_spimaster1_ointerface1_data0;
assign main_spimaster1_ointerface1_busy0 = (~main_spimaster1_spimachine1_writable0);
assign main_spimaster1_iinterface1_stb0 = (main_spimaster1_spimachine1_readable0 & main_spimaster1_read0);
assign main_spimaster1_iinterface1_data0 = main_spimaster1_spimachine1_pdi0;
assign main_spimaster1_interface_sdi0 = (main_spimaster1_interface_half_duplex0 ? main_spimaster1_interface_mosi_reg0 : main_spimaster1_interface_miso_reg0);
assign main_spimaster1_spimachine1_ce0 = (main_spimaster1_spimachine1_done0 & main_spimaster1_spimachine1_count0);
assign main_spimaster1_spimachine1_pdi0 = (main_spimaster1_spimachine1_lsb_first0 ? {main_spimaster1_spimachine1_sdi0, main_spimaster1_spimachine1_sr0[31:1]} : {main_spimaster1_spimachine1_sr0[30:0], main_spimaster1_spimachine1_sdi0});
assign main_spimaster1_spimachine1_cnt_done0 = (main_spimaster1_spimachine1_cnt0 == 1'd0);
assign main_spimaster1_spimachine1_done0 = (main_spimaster1_spimachine1_cnt_done0 & (~main_spimaster1_spimachine1_do_extend0));

// synthesis translate_off
reg dummy_d_86;
// synthesis translate_on
always @(*) begin
	main_spimaster1_spimachine1_clk_next0 <= 1'd0;
	main_spimaster1_spimachine1_cs_next0 <= 1'd0;
	main_spimaster1_spimachine1_idle0 <= 1'd0;
	main_spimaster1_spimachine1_readable0 <= 1'd0;
	main_spimaster1_spimachine1_writable0 <= 1'd0;
	main_spimaster1_spimachine1_load1 <= 1'd0;
	main_spimaster1_spimachine1_shift0 <= 1'd0;
	main_spimaster1_spimachine1_sample0 <= 1'd0;
	main_spimaster1_spimachine1_extend0 <= 1'd0;
	main_spimaster1_spimachine1_count0 <= 1'd0;
	builder_spimaster1_next_state <= 3'd0;
	builder_spimaster1_next_state <= builder_spimaster1_state;
	case (builder_spimaster1_state)
		1'd1: begin
			main_spimaster1_spimachine1_cs_next0 <= 1'd1;
			main_spimaster1_spimachine1_count0 <= 1'd1;
			main_spimaster1_spimachine1_extend0 <= 1'd1;
			main_spimaster1_spimachine1_clk_next0 <= 1'd1;
			if (main_spimaster1_spimachine1_done0) begin
				builder_spimaster1_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster1_spimachine1_cs_next0 <= 1'd1;
			main_spimaster1_spimachine1_count0 <= 1'd1;
			main_spimaster1_spimachine1_clk_next0 <= (~main_spimaster1_spimachine1_clk_phase0);
			if (main_spimaster1_spimachine1_done0) begin
				main_spimaster1_spimachine1_sample0 <= 1'd1;
				builder_spimaster1_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster1_spimachine1_cs_next0 <= 1'd1;
			main_spimaster1_spimachine1_count0 <= 1'd1;
			main_spimaster1_spimachine1_extend0 <= 1'd1;
			main_spimaster1_spimachine1_clk_next0 <= main_spimaster1_spimachine1_clk_phase0;
			if (main_spimaster1_spimachine1_done0) begin
				if ((main_spimaster1_spimachine1_n0 == 1'd0)) begin
					main_spimaster1_spimachine1_readable0 <= 1'd1;
					main_spimaster1_spimachine1_writable0 <= 1'd1;
					if (main_spimaster1_spimachine1_end1) begin
						main_spimaster1_spimachine1_clk_next0 <= 1'd0;
						main_spimaster1_spimachine1_writable0 <= 1'd0;
						if (main_spimaster1_spimachine1_clk_phase0) begin
							main_spimaster1_spimachine1_cs_next0 <= 1'd0;
							builder_spimaster1_next_state <= 3'd5;
						end else begin
							builder_spimaster1_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster1_spimachine1_load0) begin
							main_spimaster1_spimachine1_load1 <= 1'd1;
							builder_spimaster1_next_state <= 2'd2;
						end else begin
							main_spimaster1_spimachine1_count0 <= 1'd0;
						end
					end
				end else begin
					main_spimaster1_spimachine1_shift0 <= 1'd1;
					builder_spimaster1_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster1_spimachine1_count0 <= 1'd1;
			if (main_spimaster1_spimachine1_done0) begin
				builder_spimaster1_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster1_spimachine1_done0) begin
				builder_spimaster1_next_state <= 1'd0;
			end else begin
				main_spimaster1_spimachine1_count0 <= 1'd1;
			end
		end
		default: begin
			main_spimaster1_spimachine1_idle0 <= 1'd1;
			main_spimaster1_spimachine1_writable0 <= 1'd1;
			main_spimaster1_spimachine1_cs_next0 <= 1'd1;
			if (main_spimaster1_spimachine1_load0) begin
				main_spimaster1_spimachine1_count0 <= 1'd1;
				main_spimaster1_spimachine1_load1 <= 1'd1;
				if (main_spimaster1_spimachine1_clk_phase0) begin
					builder_spimaster1_next_state <= 1'd1;
				end else begin
					main_spimaster1_spimachine1_extend0 <= 1'd1;
					builder_spimaster1_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_86 <= dummy_s;
// synthesis translate_on
end
assign main_urukulmonitor1_ch_sel0 = (((main_urukulmonitor1_cs == 2'd3) | (main_urukulmonitor1_cs == 3'd4)) & (main_urukulmonitor1_current_address == 1'd0));
assign main_urukulmonitor1_ch_sel1 = (((main_urukulmonitor1_cs == 2'd3) | (main_urukulmonitor1_cs == 3'd5)) & (main_urukulmonitor1_current_address == 1'd0));
assign main_urukulmonitor1_ch_sel2 = (((main_urukulmonitor1_cs == 2'd3) | (main_urukulmonitor1_cs == 3'd6)) & (main_urukulmonitor1_current_address == 1'd0));
assign main_urukulmonitor1_ch_sel3 = (((main_urukulmonitor1_cs == 2'd3) | (main_urukulmonitor1_cs == 3'd7)) & (main_urukulmonitor1_current_address == 1'd0));

// synthesis translate_off
reg dummy_d_87;
// synthesis translate_on
always @(*) begin
	builder_ad9912monitor0_next_state <= 1'd0;
	builder_ad9912monitor0_t_next_value <= 16'd0;
	builder_ad9912monitor0_t_next_value_ce <= 1'd0;
	builder_ad9912monitor0_f_next_value <= 16'd0;
	builder_ad9912monitor0_f_next_value_ce <= 1'd0;
	builder_ad9912monitor0_next_state <= builder_ad9912monitor0_state;
	case (builder_ad9912monitor0_state)
		1'd1: begin
			if (main_urukulmonitor1_ch_sel0) begin
				if ((main_urukulmonitor1_flags & 2'd2)) begin
					builder_ad9912monitor0_t_next_value <= main_urukulmonitor1_current_data[31:16];
					builder_ad9912monitor0_t_next_value_ce <= 1'd1;
					builder_ad9912monitor0_next_state <= 1'd0;
				end else begin
					builder_ad9912monitor0_f_next_value <= main_urukulmonitor1_current_data[15:0];
					builder_ad9912monitor0_f_next_value_ce <= 1'd1;
				end
			end
		end
		default: begin
			if ((main_urukulmonitor1_ch_sel0 & (~main_urukulmonitor1_current_data[31]))) begin
				if (((main_urukulmonitor1_data_length == 5'd16) & (main_urukulmonitor1_current_data[28:16] == 9'd429))) begin
					builder_ad9912monitor0_next_state <= 1'd1;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_87 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_88;
// synthesis translate_on
always @(*) begin
	builder_ad9912monitor1_next_state <= 1'd0;
	builder_ad9912monitor1_t_next_value <= 16'd0;
	builder_ad9912monitor1_t_next_value_ce <= 1'd0;
	builder_ad9912monitor1_f_next_value <= 16'd0;
	builder_ad9912monitor1_f_next_value_ce <= 1'd0;
	builder_ad9912monitor1_next_state <= builder_ad9912monitor1_state;
	case (builder_ad9912monitor1_state)
		1'd1: begin
			if (main_urukulmonitor1_ch_sel1) begin
				if ((main_urukulmonitor1_flags & 2'd2)) begin
					builder_ad9912monitor1_t_next_value <= main_urukulmonitor1_current_data[31:16];
					builder_ad9912monitor1_t_next_value_ce <= 1'd1;
					builder_ad9912monitor1_next_state <= 1'd0;
				end else begin
					builder_ad9912monitor1_f_next_value <= main_urukulmonitor1_current_data[15:0];
					builder_ad9912monitor1_f_next_value_ce <= 1'd1;
				end
			end
		end
		default: begin
			if ((main_urukulmonitor1_ch_sel1 & (~main_urukulmonitor1_current_data[31]))) begin
				if (((main_urukulmonitor1_data_length == 5'd16) & (main_urukulmonitor1_current_data[28:16] == 9'd429))) begin
					builder_ad9912monitor1_next_state <= 1'd1;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_88 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_89;
// synthesis translate_on
always @(*) begin
	builder_ad9912monitor2_next_state <= 1'd0;
	builder_ad9912monitor2_t_next_value <= 16'd0;
	builder_ad9912monitor2_t_next_value_ce <= 1'd0;
	builder_ad9912monitor2_f_next_value <= 16'd0;
	builder_ad9912monitor2_f_next_value_ce <= 1'd0;
	builder_ad9912monitor2_next_state <= builder_ad9912monitor2_state;
	case (builder_ad9912monitor2_state)
		1'd1: begin
			if (main_urukulmonitor1_ch_sel2) begin
				if ((main_urukulmonitor1_flags & 2'd2)) begin
					builder_ad9912monitor2_t_next_value <= main_urukulmonitor1_current_data[31:16];
					builder_ad9912monitor2_t_next_value_ce <= 1'd1;
					builder_ad9912monitor2_next_state <= 1'd0;
				end else begin
					builder_ad9912monitor2_f_next_value <= main_urukulmonitor1_current_data[15:0];
					builder_ad9912monitor2_f_next_value_ce <= 1'd1;
				end
			end
		end
		default: begin
			if ((main_urukulmonitor1_ch_sel2 & (~main_urukulmonitor1_current_data[31]))) begin
				if (((main_urukulmonitor1_data_length == 5'd16) & (main_urukulmonitor1_current_data[28:16] == 9'd429))) begin
					builder_ad9912monitor2_next_state <= 1'd1;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_89 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_90;
// synthesis translate_on
always @(*) begin
	builder_ad9912monitor3_next_state <= 1'd0;
	builder_ad9912monitor3_t_next_value <= 16'd0;
	builder_ad9912monitor3_t_next_value_ce <= 1'd0;
	builder_ad9912monitor3_f_next_value <= 16'd0;
	builder_ad9912monitor3_f_next_value_ce <= 1'd0;
	builder_ad9912monitor3_next_state <= builder_ad9912monitor3_state;
	case (builder_ad9912monitor3_state)
		1'd1: begin
			if (main_urukulmonitor1_ch_sel3) begin
				if ((main_urukulmonitor1_flags & 2'd2)) begin
					builder_ad9912monitor3_t_next_value <= main_urukulmonitor1_current_data[31:16];
					builder_ad9912monitor3_t_next_value_ce <= 1'd1;
					builder_ad9912monitor3_next_state <= 1'd0;
				end else begin
					builder_ad9912monitor3_f_next_value <= main_urukulmonitor1_current_data[15:0];
					builder_ad9912monitor3_f_next_value_ce <= 1'd1;
				end
			end
		end
		default: begin
			if ((main_urukulmonitor1_ch_sel3 & (~main_urukulmonitor1_current_data[31]))) begin
				if (((main_urukulmonitor1_data_length == 5'd16) & (main_urukulmonitor1_current_data[28:16] == 9'd429))) begin
					builder_ad9912monitor3_next_state <= 1'd1;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_90 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster0_spimachine0_length1 = main_spimaster0_config_length1;
assign main_spimaster0_spimachine0_end2 = main_spimaster0_config_end1;
assign main_spimaster0_spimachine0_div1 = main_spimaster0_config_div1;
assign main_spimaster0_spimachine0_clk_phase1 = main_spimaster0_config_clk_phase1;
assign main_spimaster0_spimachine0_lsb_first1 = main_spimaster0_config_lsb_first1;
assign main_spimaster0_interface_half_duplex1 = main_spimaster0_config_half_duplex1;
assign main_spimaster0_interface_cs2 = main_spimaster0_config_cs1;
assign main_spimaster0_interface_cs_polarity1 = {1{main_spimaster0_config_cs_polarity1}};
assign main_spimaster0_interface_clk_polarity1 = main_spimaster0_config_clk_polarity1;
assign main_spimaster0_interface_offline1 = main_spimaster0_config_offline1;
assign main_spimaster0_interface_cs_next1 = main_spimaster0_spimachine0_cs_next1;
assign main_spimaster0_interface_clk_next1 = main_spimaster0_spimachine0_clk_next1;
assign main_spimaster0_interface_ce1 = main_spimaster0_spimachine0_ce1;
assign main_spimaster0_interface_sample1 = main_spimaster0_spimachine0_sample1;
assign main_spimaster0_spimachine0_sdi1 = main_spimaster0_interface_sdi1;
assign main_spimaster0_interface_sdo1 = main_spimaster0_spimachine0_sdo1;
assign main_spimaster0_spimachine0_load2 = ((main_spimaster0_ointerface0_stb1 & main_spimaster0_spimachine0_writable1) & (~main_spimaster0_ointerface0_address1));
assign main_spimaster0_spimachine0_pdo1 = main_spimaster0_ointerface0_data1;
assign main_spimaster0_ointerface0_busy1 = (~main_spimaster0_spimachine0_writable1);
assign main_spimaster0_iinterface0_stb1 = (main_spimaster0_spimachine0_readable1 & main_spimaster0_read1);
assign main_spimaster0_iinterface0_data1 = main_spimaster0_spimachine0_pdi1;
assign main_spimaster0_interface_sdi1 = (main_spimaster0_interface_half_duplex1 ? main_spimaster0_interface_mosi_reg1 : main_spimaster0_interface_miso_reg1);
assign main_spimaster0_spimachine0_ce1 = (main_spimaster0_spimachine0_done1 & main_spimaster0_spimachine0_count1);
assign main_spimaster0_spimachine0_pdi1 = (main_spimaster0_spimachine0_lsb_first1 ? {main_spimaster0_spimachine0_sdi1, main_spimaster0_spimachine0_sr1[31:1]} : {main_spimaster0_spimachine0_sr1[30:0], main_spimaster0_spimachine0_sdi1});
assign main_spimaster0_spimachine0_cnt_done1 = (main_spimaster0_spimachine0_cnt1 == 1'd0);
assign main_spimaster0_spimachine0_done1 = (main_spimaster0_spimachine0_cnt_done1 & (~main_spimaster0_spimachine0_do_extend1));

// synthesis translate_off
reg dummy_d_91;
// synthesis translate_on
always @(*) begin
	main_spimaster0_spimachine0_clk_next1 <= 1'd0;
	main_spimaster0_spimachine0_cs_next1 <= 1'd0;
	main_spimaster0_spimachine0_idle1 <= 1'd0;
	main_spimaster0_spimachine0_readable1 <= 1'd0;
	main_spimaster0_spimachine0_writable1 <= 1'd0;
	main_spimaster0_spimachine0_load3 <= 1'd0;
	main_spimaster0_spimachine0_shift1 <= 1'd0;
	main_spimaster0_spimachine0_sample1 <= 1'd0;
	main_spimaster0_spimachine0_extend1 <= 1'd0;
	main_spimaster0_spimachine0_count1 <= 1'd0;
	builder_spimaster2_next_state <= 3'd0;
	builder_spimaster2_next_state <= builder_spimaster2_state;
	case (builder_spimaster2_state)
		1'd1: begin
			main_spimaster0_spimachine0_cs_next1 <= 1'd1;
			main_spimaster0_spimachine0_count1 <= 1'd1;
			main_spimaster0_spimachine0_extend1 <= 1'd1;
			main_spimaster0_spimachine0_clk_next1 <= 1'd1;
			if (main_spimaster0_spimachine0_done1) begin
				builder_spimaster2_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster0_spimachine0_cs_next1 <= 1'd1;
			main_spimaster0_spimachine0_count1 <= 1'd1;
			main_spimaster0_spimachine0_clk_next1 <= (~main_spimaster0_spimachine0_clk_phase1);
			if (main_spimaster0_spimachine0_done1) begin
				main_spimaster0_spimachine0_sample1 <= 1'd1;
				builder_spimaster2_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster0_spimachine0_cs_next1 <= 1'd1;
			main_spimaster0_spimachine0_count1 <= 1'd1;
			main_spimaster0_spimachine0_extend1 <= 1'd1;
			main_spimaster0_spimachine0_clk_next1 <= main_spimaster0_spimachine0_clk_phase1;
			if (main_spimaster0_spimachine0_done1) begin
				if ((main_spimaster0_spimachine0_n1 == 1'd0)) begin
					main_spimaster0_spimachine0_readable1 <= 1'd1;
					main_spimaster0_spimachine0_writable1 <= 1'd1;
					if (main_spimaster0_spimachine0_end3) begin
						main_spimaster0_spimachine0_clk_next1 <= 1'd0;
						main_spimaster0_spimachine0_writable1 <= 1'd0;
						if (main_spimaster0_spimachine0_clk_phase1) begin
							main_spimaster0_spimachine0_cs_next1 <= 1'd0;
							builder_spimaster2_next_state <= 3'd5;
						end else begin
							builder_spimaster2_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster0_spimachine0_load2) begin
							main_spimaster0_spimachine0_load3 <= 1'd1;
							builder_spimaster2_next_state <= 2'd2;
						end else begin
							main_spimaster0_spimachine0_count1 <= 1'd0;
						end
					end
				end else begin
					main_spimaster0_spimachine0_shift1 <= 1'd1;
					builder_spimaster2_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster0_spimachine0_count1 <= 1'd1;
			if (main_spimaster0_spimachine0_done1) begin
				builder_spimaster2_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster0_spimachine0_done1) begin
				builder_spimaster2_next_state <= 1'd0;
			end else begin
				main_spimaster0_spimachine0_count1 <= 1'd1;
			end
		end
		default: begin
			main_spimaster0_spimachine0_idle1 <= 1'd1;
			main_spimaster0_spimachine0_writable1 <= 1'd1;
			main_spimaster0_spimachine0_cs_next1 <= 1'd1;
			if (main_spimaster0_spimachine0_load2) begin
				main_spimaster0_spimachine0_count1 <= 1'd1;
				main_spimaster0_spimachine0_load3 <= 1'd1;
				if (main_spimaster0_spimachine0_clk_phase1) begin
					builder_spimaster2_next_state <= 1'd1;
				end else begin
					main_spimaster0_spimachine0_extend1 <= 1'd1;
					builder_spimaster2_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_91 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster1_spimachine1_length1 = main_spimaster1_config_length1;
assign main_spimaster1_spimachine1_end2 = main_spimaster1_config_end1;
assign main_spimaster1_spimachine1_div1 = main_spimaster1_config_div1;
assign main_spimaster1_spimachine1_clk_phase1 = main_spimaster1_config_clk_phase1;
assign main_spimaster1_spimachine1_lsb_first1 = main_spimaster1_config_lsb_first1;
assign main_spimaster1_interface_half_duplex1 = main_spimaster1_config_half_duplex1;
assign main_spimaster1_interface_cs2 = main_spimaster1_config_cs1;
assign main_spimaster1_interface_cs_polarity1 = {1{main_spimaster1_config_cs_polarity1}};
assign main_spimaster1_interface_clk_polarity1 = main_spimaster1_config_clk_polarity1;
assign main_spimaster1_interface_offline1 = main_spimaster1_config_offline1;
assign main_spimaster1_interface_cs_next1 = main_spimaster1_spimachine1_cs_next1;
assign main_spimaster1_interface_clk_next1 = main_spimaster1_spimachine1_clk_next1;
assign main_spimaster1_interface_ce1 = main_spimaster1_spimachine1_ce1;
assign main_spimaster1_interface_sample1 = main_spimaster1_spimachine1_sample1;
assign main_spimaster1_spimachine1_sdi1 = main_spimaster1_interface_sdi1;
assign main_spimaster1_interface_sdo1 = main_spimaster1_spimachine1_sdo1;
assign main_spimaster1_spimachine1_load2 = ((main_spimaster1_ointerface1_stb1 & main_spimaster1_spimachine1_writable1) & (~main_spimaster1_ointerface1_address1));
assign main_spimaster1_spimachine1_pdo1 = main_spimaster1_ointerface1_data1;
assign main_spimaster1_ointerface1_busy1 = (~main_spimaster1_spimachine1_writable1);
assign main_spimaster1_iinterface1_stb1 = (main_spimaster1_spimachine1_readable1 & main_spimaster1_read1);
assign main_spimaster1_iinterface1_data1 = main_spimaster1_spimachine1_pdi1;
assign main_spimaster1_interface_sdi1 = (main_spimaster1_interface_half_duplex1 ? main_spimaster1_interface_mosi_reg1 : main_spimaster1_interface_miso_reg1);
assign main_spimaster1_spimachine1_ce1 = (main_spimaster1_spimachine1_done1 & main_spimaster1_spimachine1_count1);
assign main_spimaster1_spimachine1_pdi1 = (main_spimaster1_spimachine1_lsb_first1 ? {main_spimaster1_spimachine1_sdi1, main_spimaster1_spimachine1_sr1[31:1]} : {main_spimaster1_spimachine1_sr1[30:0], main_spimaster1_spimachine1_sdi1});
assign main_spimaster1_spimachine1_cnt_done1 = (main_spimaster1_spimachine1_cnt1 == 1'd0);
assign main_spimaster1_spimachine1_done1 = (main_spimaster1_spimachine1_cnt_done1 & (~main_spimaster1_spimachine1_do_extend1));

// synthesis translate_off
reg dummy_d_92;
// synthesis translate_on
always @(*) begin
	main_spimaster1_spimachine1_clk_next1 <= 1'd0;
	main_spimaster1_spimachine1_cs_next1 <= 1'd0;
	main_spimaster1_spimachine1_idle1 <= 1'd0;
	main_spimaster1_spimachine1_readable1 <= 1'd0;
	main_spimaster1_spimachine1_writable1 <= 1'd0;
	main_spimaster1_spimachine1_load3 <= 1'd0;
	main_spimaster1_spimachine1_shift1 <= 1'd0;
	main_spimaster1_spimachine1_sample1 <= 1'd0;
	main_spimaster1_spimachine1_extend1 <= 1'd0;
	main_spimaster1_spimachine1_count1 <= 1'd0;
	builder_spimaster3_next_state <= 3'd0;
	builder_spimaster3_next_state <= builder_spimaster3_state;
	case (builder_spimaster3_state)
		1'd1: begin
			main_spimaster1_spimachine1_cs_next1 <= 1'd1;
			main_spimaster1_spimachine1_count1 <= 1'd1;
			main_spimaster1_spimachine1_extend1 <= 1'd1;
			main_spimaster1_spimachine1_clk_next1 <= 1'd1;
			if (main_spimaster1_spimachine1_done1) begin
				builder_spimaster3_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster1_spimachine1_cs_next1 <= 1'd1;
			main_spimaster1_spimachine1_count1 <= 1'd1;
			main_spimaster1_spimachine1_clk_next1 <= (~main_spimaster1_spimachine1_clk_phase1);
			if (main_spimaster1_spimachine1_done1) begin
				main_spimaster1_spimachine1_sample1 <= 1'd1;
				builder_spimaster3_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster1_spimachine1_cs_next1 <= 1'd1;
			main_spimaster1_spimachine1_count1 <= 1'd1;
			main_spimaster1_spimachine1_extend1 <= 1'd1;
			main_spimaster1_spimachine1_clk_next1 <= main_spimaster1_spimachine1_clk_phase1;
			if (main_spimaster1_spimachine1_done1) begin
				if ((main_spimaster1_spimachine1_n1 == 1'd0)) begin
					main_spimaster1_spimachine1_readable1 <= 1'd1;
					main_spimaster1_spimachine1_writable1 <= 1'd1;
					if (main_spimaster1_spimachine1_end3) begin
						main_spimaster1_spimachine1_clk_next1 <= 1'd0;
						main_spimaster1_spimachine1_writable1 <= 1'd0;
						if (main_spimaster1_spimachine1_clk_phase1) begin
							main_spimaster1_spimachine1_cs_next1 <= 1'd0;
							builder_spimaster3_next_state <= 3'd5;
						end else begin
							builder_spimaster3_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster1_spimachine1_load2) begin
							main_spimaster1_spimachine1_load3 <= 1'd1;
							builder_spimaster3_next_state <= 2'd2;
						end else begin
							main_spimaster1_spimachine1_count1 <= 1'd0;
						end
					end
				end else begin
					main_spimaster1_spimachine1_shift1 <= 1'd1;
					builder_spimaster3_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster1_spimachine1_count1 <= 1'd1;
			if (main_spimaster1_spimachine1_done1) begin
				builder_spimaster3_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster1_spimachine1_done1) begin
				builder_spimaster3_next_state <= 1'd0;
			end else begin
				main_spimaster1_spimachine1_count1 <= 1'd1;
			end
		end
		default: begin
			main_spimaster1_spimachine1_idle1 <= 1'd1;
			main_spimaster1_spimachine1_writable1 <= 1'd1;
			main_spimaster1_spimachine1_cs_next1 <= 1'd1;
			if (main_spimaster1_spimachine1_load2) begin
				main_spimaster1_spimachine1_count1 <= 1'd1;
				main_spimaster1_spimachine1_load3 <= 1'd1;
				if (main_spimaster1_spimachine1_clk_phase1) begin
					builder_spimaster3_next_state <= 1'd1;
				end else begin
					main_spimaster1_spimachine1_extend1 <= 1'd1;
					builder_spimaster3_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_92 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster2_spimachine2_length = main_spimaster2_config_length;
assign main_spimaster2_spimachine2_end0 = main_spimaster2_config_end;
assign main_spimaster2_spimachine2_div = main_spimaster2_config_div;
assign main_spimaster2_spimachine2_clk_phase = main_spimaster2_config_clk_phase;
assign main_spimaster2_spimachine2_lsb_first = main_spimaster2_config_lsb_first;
assign main_spimaster2_interface_half_duplex = main_spimaster2_config_half_duplex;
assign main_spimaster2_interface_cs0 = main_spimaster2_config_cs;
assign main_spimaster2_interface_cs_polarity = {2{main_spimaster2_config_cs_polarity}};
assign main_spimaster2_interface_clk_polarity = main_spimaster2_config_clk_polarity;
assign main_spimaster2_interface_offline = main_spimaster2_config_offline;
assign main_spimaster2_interface_cs_next = main_spimaster2_spimachine2_cs_next;
assign main_spimaster2_interface_clk_next = main_spimaster2_spimachine2_clk_next;
assign main_spimaster2_interface_ce = main_spimaster2_spimachine2_ce;
assign main_spimaster2_interface_sample = main_spimaster2_spimachine2_sample;
assign main_spimaster2_spimachine2_sdi = main_spimaster2_interface_sdi;
assign main_spimaster2_interface_sdo = main_spimaster2_spimachine2_sdo;
assign main_spimaster2_spimachine2_load0 = ((main_spimaster2_ointerface2_stb & main_spimaster2_spimachine2_writable) & (~main_spimaster2_ointerface2_address));
assign main_spimaster2_spimachine2_pdo = main_spimaster2_ointerface2_data;
assign main_spimaster2_ointerface2_busy = (~main_spimaster2_spimachine2_writable);
assign main_spimaster2_iinterface2_stb = (main_spimaster2_spimachine2_readable & main_spimaster2_read);
assign main_spimaster2_iinterface2_data = main_spimaster2_spimachine2_pdi;
assign main_spimaster2_interface_sdi = (main_spimaster2_interface_half_duplex ? main_spimaster2_interface_mosi_reg : main_spimaster2_interface_miso_reg);
assign main_spimaster2_spimachine2_ce = (main_spimaster2_spimachine2_done & main_spimaster2_spimachine2_count);
assign main_spimaster2_spimachine2_pdi = (main_spimaster2_spimachine2_lsb_first ? {main_spimaster2_spimachine2_sdi, main_spimaster2_spimachine2_sr[31:1]} : {main_spimaster2_spimachine2_sr[30:0], main_spimaster2_spimachine2_sdi});
assign main_spimaster2_spimachine2_cnt_done = (main_spimaster2_spimachine2_cnt == 1'd0);
assign main_spimaster2_spimachine2_done = (main_spimaster2_spimachine2_cnt_done & (~main_spimaster2_spimachine2_do_extend));

// synthesis translate_off
reg dummy_d_93;
// synthesis translate_on
always @(*) begin
	main_spimaster2_spimachine2_clk_next <= 1'd0;
	main_spimaster2_spimachine2_cs_next <= 1'd0;
	main_spimaster2_spimachine2_idle <= 1'd0;
	main_spimaster2_spimachine2_readable <= 1'd0;
	main_spimaster2_spimachine2_writable <= 1'd0;
	main_spimaster2_spimachine2_load1 <= 1'd0;
	main_spimaster2_spimachine2_shift <= 1'd0;
	main_spimaster2_spimachine2_sample <= 1'd0;
	main_spimaster2_spimachine2_extend <= 1'd0;
	main_spimaster2_spimachine2_count <= 1'd0;
	builder_spimaster4_next_state <= 3'd0;
	builder_spimaster4_next_state <= builder_spimaster4_state;
	case (builder_spimaster4_state)
		1'd1: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_extend <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= 1'd1;
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster4_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= (~main_spimaster2_spimachine2_clk_phase);
			if (main_spimaster2_spimachine2_done) begin
				main_spimaster2_spimachine2_sample <= 1'd1;
				builder_spimaster4_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_extend <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= main_spimaster2_spimachine2_clk_phase;
			if (main_spimaster2_spimachine2_done) begin
				if ((main_spimaster2_spimachine2_n == 1'd0)) begin
					main_spimaster2_spimachine2_readable <= 1'd1;
					main_spimaster2_spimachine2_writable <= 1'd1;
					if (main_spimaster2_spimachine2_end1) begin
						main_spimaster2_spimachine2_clk_next <= 1'd0;
						main_spimaster2_spimachine2_writable <= 1'd0;
						if (main_spimaster2_spimachine2_clk_phase) begin
							main_spimaster2_spimachine2_cs_next <= 1'd0;
							builder_spimaster4_next_state <= 3'd5;
						end else begin
							builder_spimaster4_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster2_spimachine2_load0) begin
							main_spimaster2_spimachine2_load1 <= 1'd1;
							builder_spimaster4_next_state <= 2'd2;
						end else begin
							main_spimaster2_spimachine2_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster2_spimachine2_shift <= 1'd1;
					builder_spimaster4_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster2_spimachine2_count <= 1'd1;
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster4_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster4_next_state <= 1'd0;
			end else begin
				main_spimaster2_spimachine2_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster2_spimachine2_idle <= 1'd1;
			main_spimaster2_spimachine2_writable <= 1'd1;
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			if (main_spimaster2_spimachine2_load0) begin
				main_spimaster2_spimachine2_count <= 1'd1;
				main_spimaster2_spimachine2_load1 <= 1'd1;
				if (main_spimaster2_spimachine2_clk_phase) begin
					builder_spimaster4_next_state <= 1'd1;
				end else begin
					main_spimaster2_spimachine2_extend <= 1'd1;
					builder_spimaster4_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_93 <= dummy_s;
// synthesis translate_on
end
assign user_led = main_output0_pad_o;
assign user_led_1 = main_output1_pad_o;
assign user_led_2 = main_output2_pad_o;
assign main_genericstandalone_full_ts = (main_genericstandalone_coarse_ts <<< 2'd3);
assign rio_clk = sys_clk;
assign rio_rst = main_genericstandalone_rtio_core_cmd_reset;
assign rio_phy_clk = sys_clk;
assign rio_phy_rst = main_genericstandalone_rtio_core_cmd_reset_phy;
assign main_genericstandalone_rtio_core_sed_gates_coarse_timestamp = main_genericstandalone_coarse_ts;
assign main_genericstandalone_rtio_core_async_error_w = {main_genericstandalone_rtio_core_o_sequence_error, main_genericstandalone_rtio_core_o_busy, main_genericstandalone_rtio_core_o_collision};
assign main_genericstandalone_rtio_core_o_collision_sync_i = main_genericstandalone_rtio_core_sed_collision;
assign main_genericstandalone_rtio_core_o_collision_sync_data_i = main_genericstandalone_rtio_core_sed_collision_channel;
assign main_genericstandalone_rtio_core_o_busy_sync_i = main_genericstandalone_rtio_core_sed_busy;
assign main_genericstandalone_rtio_core_o_busy_sync_data_i = main_genericstandalone_rtio_core_sed_busy_channel;
assign main_genericstandalone_rtio_core_sed_record0_we = main_genericstandalone_rtio_core_sed_lane_dist_record0_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record0_writable = main_genericstandalone_rtio_core_sed_record0_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record0_high_watermark = main_genericstandalone_rtio_core_sed_record0_high_watermark;
assign main_genericstandalone_rtio_core_sed_record0_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record0_seqn;
assign main_genericstandalone_rtio_core_sed_record0_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_channel;
assign main_genericstandalone_rtio_core_sed_record0_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record0_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_address;
assign main_genericstandalone_rtio_core_sed_record0_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_data;
assign main_genericstandalone_rtio_core_sed_record1_we = main_genericstandalone_rtio_core_sed_lane_dist_record1_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record1_writable = main_genericstandalone_rtio_core_sed_record1_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record1_high_watermark = main_genericstandalone_rtio_core_sed_record1_high_watermark;
assign main_genericstandalone_rtio_core_sed_record1_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record1_seqn;
assign main_genericstandalone_rtio_core_sed_record1_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_channel;
assign main_genericstandalone_rtio_core_sed_record1_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record1_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_address;
assign main_genericstandalone_rtio_core_sed_record1_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_data;
assign main_genericstandalone_rtio_core_sed_record2_we = main_genericstandalone_rtio_core_sed_lane_dist_record2_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record2_writable = main_genericstandalone_rtio_core_sed_record2_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record2_high_watermark = main_genericstandalone_rtio_core_sed_record2_high_watermark;
assign main_genericstandalone_rtio_core_sed_record2_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record2_seqn;
assign main_genericstandalone_rtio_core_sed_record2_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_channel;
assign main_genericstandalone_rtio_core_sed_record2_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record2_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_address;
assign main_genericstandalone_rtio_core_sed_record2_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_data;
assign main_genericstandalone_rtio_core_sed_record3_we = main_genericstandalone_rtio_core_sed_lane_dist_record3_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record3_writable = main_genericstandalone_rtio_core_sed_record3_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record3_high_watermark = main_genericstandalone_rtio_core_sed_record3_high_watermark;
assign main_genericstandalone_rtio_core_sed_record3_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record3_seqn;
assign main_genericstandalone_rtio_core_sed_record3_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_channel;
assign main_genericstandalone_rtio_core_sed_record3_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record3_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_address;
assign main_genericstandalone_rtio_core_sed_record3_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_data;
assign main_genericstandalone_rtio_core_sed_record4_we = main_genericstandalone_rtio_core_sed_lane_dist_record4_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record4_writable = main_genericstandalone_rtio_core_sed_record4_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record4_high_watermark = main_genericstandalone_rtio_core_sed_record4_high_watermark;
assign main_genericstandalone_rtio_core_sed_record4_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record4_seqn;
assign main_genericstandalone_rtio_core_sed_record4_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_channel;
assign main_genericstandalone_rtio_core_sed_record4_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record4_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_address;
assign main_genericstandalone_rtio_core_sed_record4_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_data;
assign main_genericstandalone_rtio_core_sed_record5_we = main_genericstandalone_rtio_core_sed_lane_dist_record5_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record5_writable = main_genericstandalone_rtio_core_sed_record5_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record5_high_watermark = main_genericstandalone_rtio_core_sed_record5_high_watermark;
assign main_genericstandalone_rtio_core_sed_record5_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record5_seqn;
assign main_genericstandalone_rtio_core_sed_record5_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_channel;
assign main_genericstandalone_rtio_core_sed_record5_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record5_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_address;
assign main_genericstandalone_rtio_core_sed_record5_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_data;
assign main_genericstandalone_rtio_core_sed_record6_we = main_genericstandalone_rtio_core_sed_lane_dist_record6_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record6_writable = main_genericstandalone_rtio_core_sed_record6_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record6_high_watermark = main_genericstandalone_rtio_core_sed_record6_high_watermark;
assign main_genericstandalone_rtio_core_sed_record6_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record6_seqn;
assign main_genericstandalone_rtio_core_sed_record6_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_channel;
assign main_genericstandalone_rtio_core_sed_record6_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record6_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_address;
assign main_genericstandalone_rtio_core_sed_record6_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_data;
assign main_genericstandalone_rtio_core_sed_record7_we = main_genericstandalone_rtio_core_sed_lane_dist_record7_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record7_writable = main_genericstandalone_rtio_core_sed_record7_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record7_high_watermark = main_genericstandalone_rtio_core_sed_record7_high_watermark;
assign main_genericstandalone_rtio_core_sed_record7_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record7_seqn;
assign main_genericstandalone_rtio_core_sed_record7_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_channel;
assign main_genericstandalone_rtio_core_sed_record7_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record7_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_address;
assign main_genericstandalone_rtio_core_sed_record7_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_data;
assign main_genericstandalone_rtio_core_sed_record8_we = main_genericstandalone_rtio_core_sed_lane_dist_record8_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record8_writable = main_genericstandalone_rtio_core_sed_record8_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record8_high_watermark = main_genericstandalone_rtio_core_sed_record8_high_watermark;
assign main_genericstandalone_rtio_core_sed_record8_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record8_seqn;
assign main_genericstandalone_rtio_core_sed_record8_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_channel;
assign main_genericstandalone_rtio_core_sed_record8_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record8_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_address;
assign main_genericstandalone_rtio_core_sed_record8_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_data;
assign main_genericstandalone_rtio_core_sed_record9_we = main_genericstandalone_rtio_core_sed_lane_dist_record9_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record9_writable = main_genericstandalone_rtio_core_sed_record9_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record9_high_watermark = main_genericstandalone_rtio_core_sed_record9_high_watermark;
assign main_genericstandalone_rtio_core_sed_record9_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record9_seqn;
assign main_genericstandalone_rtio_core_sed_record9_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_channel;
assign main_genericstandalone_rtio_core_sed_record9_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record9_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_address;
assign main_genericstandalone_rtio_core_sed_record9_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_data;
assign main_genericstandalone_rtio_core_sed_record10_we = main_genericstandalone_rtio_core_sed_lane_dist_record10_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record10_writable = main_genericstandalone_rtio_core_sed_record10_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record10_high_watermark = main_genericstandalone_rtio_core_sed_record10_high_watermark;
assign main_genericstandalone_rtio_core_sed_record10_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record10_seqn;
assign main_genericstandalone_rtio_core_sed_record10_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_channel;
assign main_genericstandalone_rtio_core_sed_record10_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record10_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_address;
assign main_genericstandalone_rtio_core_sed_record10_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_data;
assign main_genericstandalone_rtio_core_sed_record11_we = main_genericstandalone_rtio_core_sed_lane_dist_record11_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record11_writable = main_genericstandalone_rtio_core_sed_record11_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record11_high_watermark = main_genericstandalone_rtio_core_sed_record11_high_watermark;
assign main_genericstandalone_rtio_core_sed_record11_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record11_seqn;
assign main_genericstandalone_rtio_core_sed_record11_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_channel;
assign main_genericstandalone_rtio_core_sed_record11_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record11_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_address;
assign main_genericstandalone_rtio_core_sed_record11_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_data;
assign main_genericstandalone_rtio_core_sed_record12_we = main_genericstandalone_rtio_core_sed_lane_dist_record12_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record12_writable = main_genericstandalone_rtio_core_sed_record12_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record12_high_watermark = main_genericstandalone_rtio_core_sed_record12_high_watermark;
assign main_genericstandalone_rtio_core_sed_record12_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record12_seqn;
assign main_genericstandalone_rtio_core_sed_record12_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_channel;
assign main_genericstandalone_rtio_core_sed_record12_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record12_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_address;
assign main_genericstandalone_rtio_core_sed_record12_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_data;
assign main_genericstandalone_rtio_core_sed_record13_we = main_genericstandalone_rtio_core_sed_lane_dist_record13_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record13_writable = main_genericstandalone_rtio_core_sed_record13_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record13_high_watermark = main_genericstandalone_rtio_core_sed_record13_high_watermark;
assign main_genericstandalone_rtio_core_sed_record13_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record13_seqn;
assign main_genericstandalone_rtio_core_sed_record13_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_channel;
assign main_genericstandalone_rtio_core_sed_record13_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record13_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_address;
assign main_genericstandalone_rtio_core_sed_record13_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_data;
assign main_genericstandalone_rtio_core_sed_record14_we = main_genericstandalone_rtio_core_sed_lane_dist_record14_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record14_writable = main_genericstandalone_rtio_core_sed_record14_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record14_high_watermark = main_genericstandalone_rtio_core_sed_record14_high_watermark;
assign main_genericstandalone_rtio_core_sed_record14_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record14_seqn;
assign main_genericstandalone_rtio_core_sed_record14_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_channel;
assign main_genericstandalone_rtio_core_sed_record14_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record14_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_address;
assign main_genericstandalone_rtio_core_sed_record14_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_data;
assign main_genericstandalone_rtio_core_sed_record15_we = main_genericstandalone_rtio_core_sed_lane_dist_record15_we;
assign main_genericstandalone_rtio_core_sed_lane_dist_record15_writable = main_genericstandalone_rtio_core_sed_record15_writable;
assign main_genericstandalone_rtio_core_sed_lane_dist_record15_high_watermark = main_genericstandalone_rtio_core_sed_record15_high_watermark;
assign main_genericstandalone_rtio_core_sed_record15_seqn0 = main_genericstandalone_rtio_core_sed_lane_dist_record15_seqn;
assign main_genericstandalone_rtio_core_sed_record15_payload_channel0 = main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_channel;
assign main_genericstandalone_rtio_core_sed_record15_payload_timestamp = main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_record15_payload_address0 = main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_address;
assign main_genericstandalone_rtio_core_sed_record15_payload_data0 = main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_data;
assign main_genericstandalone_rtio_core_sed_record16_re = main_genericstandalone_rtio_core_sed_gates_record0_re;
assign main_genericstandalone_rtio_core_sed_gates_record0_readable = main_genericstandalone_rtio_core_sed_record16_readable;
assign main_genericstandalone_rtio_core_sed_gates_record0_seqn = main_genericstandalone_rtio_core_sed_record16_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record0_payload_channel = main_genericstandalone_rtio_core_sed_record16_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record0_payload_timestamp = main_genericstandalone_rtio_core_sed_record16_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record0_payload_address = main_genericstandalone_rtio_core_sed_record16_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record0_payload_data = main_genericstandalone_rtio_core_sed_record16_payload_data;
assign main_genericstandalone_rtio_core_sed_record17_re = main_genericstandalone_rtio_core_sed_gates_record1_re;
assign main_genericstandalone_rtio_core_sed_gates_record1_readable = main_genericstandalone_rtio_core_sed_record17_readable;
assign main_genericstandalone_rtio_core_sed_gates_record1_seqn = main_genericstandalone_rtio_core_sed_record17_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record1_payload_channel = main_genericstandalone_rtio_core_sed_record17_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record1_payload_timestamp = main_genericstandalone_rtio_core_sed_record17_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record1_payload_address = main_genericstandalone_rtio_core_sed_record17_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record1_payload_data = main_genericstandalone_rtio_core_sed_record17_payload_data;
assign main_genericstandalone_rtio_core_sed_record18_re = main_genericstandalone_rtio_core_sed_gates_record2_re;
assign main_genericstandalone_rtio_core_sed_gates_record2_readable = main_genericstandalone_rtio_core_sed_record18_readable;
assign main_genericstandalone_rtio_core_sed_gates_record2_seqn = main_genericstandalone_rtio_core_sed_record18_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record2_payload_channel = main_genericstandalone_rtio_core_sed_record18_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record2_payload_timestamp = main_genericstandalone_rtio_core_sed_record18_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record2_payload_address = main_genericstandalone_rtio_core_sed_record18_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record2_payload_data = main_genericstandalone_rtio_core_sed_record18_payload_data;
assign main_genericstandalone_rtio_core_sed_record19_re = main_genericstandalone_rtio_core_sed_gates_record3_re;
assign main_genericstandalone_rtio_core_sed_gates_record3_readable = main_genericstandalone_rtio_core_sed_record19_readable;
assign main_genericstandalone_rtio_core_sed_gates_record3_seqn = main_genericstandalone_rtio_core_sed_record19_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record3_payload_channel = main_genericstandalone_rtio_core_sed_record19_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record3_payload_timestamp = main_genericstandalone_rtio_core_sed_record19_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record3_payload_address = main_genericstandalone_rtio_core_sed_record19_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record3_payload_data = main_genericstandalone_rtio_core_sed_record19_payload_data;
assign main_genericstandalone_rtio_core_sed_record20_re = main_genericstandalone_rtio_core_sed_gates_record4_re;
assign main_genericstandalone_rtio_core_sed_gates_record4_readable = main_genericstandalone_rtio_core_sed_record20_readable;
assign main_genericstandalone_rtio_core_sed_gates_record4_seqn = main_genericstandalone_rtio_core_sed_record20_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record4_payload_channel = main_genericstandalone_rtio_core_sed_record20_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record4_payload_timestamp = main_genericstandalone_rtio_core_sed_record20_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record4_payload_address = main_genericstandalone_rtio_core_sed_record20_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record4_payload_data = main_genericstandalone_rtio_core_sed_record20_payload_data;
assign main_genericstandalone_rtio_core_sed_record21_re = main_genericstandalone_rtio_core_sed_gates_record5_re;
assign main_genericstandalone_rtio_core_sed_gates_record5_readable = main_genericstandalone_rtio_core_sed_record21_readable;
assign main_genericstandalone_rtio_core_sed_gates_record5_seqn = main_genericstandalone_rtio_core_sed_record21_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record5_payload_channel = main_genericstandalone_rtio_core_sed_record21_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record5_payload_timestamp = main_genericstandalone_rtio_core_sed_record21_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record5_payload_address = main_genericstandalone_rtio_core_sed_record21_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record5_payload_data = main_genericstandalone_rtio_core_sed_record21_payload_data;
assign main_genericstandalone_rtio_core_sed_record22_re = main_genericstandalone_rtio_core_sed_gates_record6_re;
assign main_genericstandalone_rtio_core_sed_gates_record6_readable = main_genericstandalone_rtio_core_sed_record22_readable;
assign main_genericstandalone_rtio_core_sed_gates_record6_seqn = main_genericstandalone_rtio_core_sed_record22_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record6_payload_channel = main_genericstandalone_rtio_core_sed_record22_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record6_payload_timestamp = main_genericstandalone_rtio_core_sed_record22_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record6_payload_address = main_genericstandalone_rtio_core_sed_record22_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record6_payload_data = main_genericstandalone_rtio_core_sed_record22_payload_data;
assign main_genericstandalone_rtio_core_sed_record23_re = main_genericstandalone_rtio_core_sed_gates_record7_re;
assign main_genericstandalone_rtio_core_sed_gates_record7_readable = main_genericstandalone_rtio_core_sed_record23_readable;
assign main_genericstandalone_rtio_core_sed_gates_record7_seqn = main_genericstandalone_rtio_core_sed_record23_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record7_payload_channel = main_genericstandalone_rtio_core_sed_record23_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record7_payload_timestamp = main_genericstandalone_rtio_core_sed_record23_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record7_payload_address = main_genericstandalone_rtio_core_sed_record23_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record7_payload_data = main_genericstandalone_rtio_core_sed_record23_payload_data;
assign main_genericstandalone_rtio_core_sed_record24_re = main_genericstandalone_rtio_core_sed_gates_record8_re;
assign main_genericstandalone_rtio_core_sed_gates_record8_readable = main_genericstandalone_rtio_core_sed_record24_readable;
assign main_genericstandalone_rtio_core_sed_gates_record8_seqn = main_genericstandalone_rtio_core_sed_record24_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record8_payload_channel = main_genericstandalone_rtio_core_sed_record24_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record8_payload_timestamp = main_genericstandalone_rtio_core_sed_record24_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record8_payload_address = main_genericstandalone_rtio_core_sed_record24_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record8_payload_data = main_genericstandalone_rtio_core_sed_record24_payload_data;
assign main_genericstandalone_rtio_core_sed_record25_re = main_genericstandalone_rtio_core_sed_gates_record9_re;
assign main_genericstandalone_rtio_core_sed_gates_record9_readable = main_genericstandalone_rtio_core_sed_record25_readable;
assign main_genericstandalone_rtio_core_sed_gates_record9_seqn = main_genericstandalone_rtio_core_sed_record25_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record9_payload_channel = main_genericstandalone_rtio_core_sed_record25_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record9_payload_timestamp = main_genericstandalone_rtio_core_sed_record25_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record9_payload_address = main_genericstandalone_rtio_core_sed_record25_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record9_payload_data = main_genericstandalone_rtio_core_sed_record25_payload_data;
assign main_genericstandalone_rtio_core_sed_record26_re = main_genericstandalone_rtio_core_sed_gates_record10_re;
assign main_genericstandalone_rtio_core_sed_gates_record10_readable = main_genericstandalone_rtio_core_sed_record26_readable;
assign main_genericstandalone_rtio_core_sed_gates_record10_seqn = main_genericstandalone_rtio_core_sed_record26_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record10_payload_channel = main_genericstandalone_rtio_core_sed_record26_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record10_payload_timestamp = main_genericstandalone_rtio_core_sed_record26_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record10_payload_address = main_genericstandalone_rtio_core_sed_record26_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record10_payload_data = main_genericstandalone_rtio_core_sed_record26_payload_data;
assign main_genericstandalone_rtio_core_sed_record27_re = main_genericstandalone_rtio_core_sed_gates_record11_re;
assign main_genericstandalone_rtio_core_sed_gates_record11_readable = main_genericstandalone_rtio_core_sed_record27_readable;
assign main_genericstandalone_rtio_core_sed_gates_record11_seqn = main_genericstandalone_rtio_core_sed_record27_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record11_payload_channel = main_genericstandalone_rtio_core_sed_record27_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record11_payload_timestamp = main_genericstandalone_rtio_core_sed_record27_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record11_payload_address = main_genericstandalone_rtio_core_sed_record27_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record11_payload_data = main_genericstandalone_rtio_core_sed_record27_payload_data;
assign main_genericstandalone_rtio_core_sed_record28_re = main_genericstandalone_rtio_core_sed_gates_record12_re;
assign main_genericstandalone_rtio_core_sed_gates_record12_readable = main_genericstandalone_rtio_core_sed_record28_readable;
assign main_genericstandalone_rtio_core_sed_gates_record12_seqn = main_genericstandalone_rtio_core_sed_record28_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record12_payload_channel = main_genericstandalone_rtio_core_sed_record28_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record12_payload_timestamp = main_genericstandalone_rtio_core_sed_record28_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record12_payload_address = main_genericstandalone_rtio_core_sed_record28_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record12_payload_data = main_genericstandalone_rtio_core_sed_record28_payload_data;
assign main_genericstandalone_rtio_core_sed_record29_re = main_genericstandalone_rtio_core_sed_gates_record13_re;
assign main_genericstandalone_rtio_core_sed_gates_record13_readable = main_genericstandalone_rtio_core_sed_record29_readable;
assign main_genericstandalone_rtio_core_sed_gates_record13_seqn = main_genericstandalone_rtio_core_sed_record29_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record13_payload_channel = main_genericstandalone_rtio_core_sed_record29_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record13_payload_timestamp = main_genericstandalone_rtio_core_sed_record29_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record13_payload_address = main_genericstandalone_rtio_core_sed_record29_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record13_payload_data = main_genericstandalone_rtio_core_sed_record29_payload_data;
assign main_genericstandalone_rtio_core_sed_record30_re = main_genericstandalone_rtio_core_sed_gates_record14_re;
assign main_genericstandalone_rtio_core_sed_gates_record14_readable = main_genericstandalone_rtio_core_sed_record30_readable;
assign main_genericstandalone_rtio_core_sed_gates_record14_seqn = main_genericstandalone_rtio_core_sed_record30_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record14_payload_channel = main_genericstandalone_rtio_core_sed_record30_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record14_payload_timestamp = main_genericstandalone_rtio_core_sed_record30_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record14_payload_address = main_genericstandalone_rtio_core_sed_record30_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record14_payload_data = main_genericstandalone_rtio_core_sed_record30_payload_data;
assign main_genericstandalone_rtio_core_sed_record31_re = main_genericstandalone_rtio_core_sed_gates_record15_re;
assign main_genericstandalone_rtio_core_sed_gates_record15_readable = main_genericstandalone_rtio_core_sed_record31_readable;
assign main_genericstandalone_rtio_core_sed_gates_record15_seqn = main_genericstandalone_rtio_core_sed_record31_seqn;
assign main_genericstandalone_rtio_core_sed_gates_record15_payload_channel = main_genericstandalone_rtio_core_sed_record31_payload_channel;
assign main_genericstandalone_rtio_core_sed_gates_record15_payload_timestamp = main_genericstandalone_rtio_core_sed_record31_payload_timestamp;
assign main_genericstandalone_rtio_core_sed_gates_record15_payload_address = main_genericstandalone_rtio_core_sed_record31_payload_address;
assign main_genericstandalone_rtio_core_sed_gates_record15_payload_data = main_genericstandalone_rtio_core_sed_record31_payload_data;
assign main_genericstandalone_rtio_core_sed_record0_valid0 = main_genericstandalone_rtio_core_sed_gates_record16_valid;
assign main_genericstandalone_rtio_core_sed_record0_seqn1 = main_genericstandalone_rtio_core_sed_gates_record16_seqn;
assign main_genericstandalone_rtio_core_sed_record0_replace_occured = main_genericstandalone_rtio_core_sed_gates_record16_replace_occured;
assign main_genericstandalone_rtio_core_sed_record0_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record16_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record0_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record16_payload_channel;
assign main_genericstandalone_rtio_core_sed_record0_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record16_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record0_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record16_payload_address;
assign main_genericstandalone_rtio_core_sed_record0_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record16_payload_data;
assign main_genericstandalone_rtio_core_sed_record1_valid0 = main_genericstandalone_rtio_core_sed_gates_record17_valid;
assign main_genericstandalone_rtio_core_sed_record1_seqn1 = main_genericstandalone_rtio_core_sed_gates_record17_seqn;
assign main_genericstandalone_rtio_core_sed_record1_replace_occured = main_genericstandalone_rtio_core_sed_gates_record17_replace_occured;
assign main_genericstandalone_rtio_core_sed_record1_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record17_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record1_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record17_payload_channel;
assign main_genericstandalone_rtio_core_sed_record1_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record17_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record1_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record17_payload_address;
assign main_genericstandalone_rtio_core_sed_record1_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record17_payload_data;
assign main_genericstandalone_rtio_core_sed_record2_valid0 = main_genericstandalone_rtio_core_sed_gates_record18_valid;
assign main_genericstandalone_rtio_core_sed_record2_seqn1 = main_genericstandalone_rtio_core_sed_gates_record18_seqn;
assign main_genericstandalone_rtio_core_sed_record2_replace_occured = main_genericstandalone_rtio_core_sed_gates_record18_replace_occured;
assign main_genericstandalone_rtio_core_sed_record2_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record18_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record2_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record18_payload_channel;
assign main_genericstandalone_rtio_core_sed_record2_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record18_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record2_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record18_payload_address;
assign main_genericstandalone_rtio_core_sed_record2_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record18_payload_data;
assign main_genericstandalone_rtio_core_sed_record3_valid0 = main_genericstandalone_rtio_core_sed_gates_record19_valid;
assign main_genericstandalone_rtio_core_sed_record3_seqn1 = main_genericstandalone_rtio_core_sed_gates_record19_seqn;
assign main_genericstandalone_rtio_core_sed_record3_replace_occured = main_genericstandalone_rtio_core_sed_gates_record19_replace_occured;
assign main_genericstandalone_rtio_core_sed_record3_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record19_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record3_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record19_payload_channel;
assign main_genericstandalone_rtio_core_sed_record3_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record19_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record3_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record19_payload_address;
assign main_genericstandalone_rtio_core_sed_record3_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record19_payload_data;
assign main_genericstandalone_rtio_core_sed_record4_valid0 = main_genericstandalone_rtio_core_sed_gates_record20_valid;
assign main_genericstandalone_rtio_core_sed_record4_seqn1 = main_genericstandalone_rtio_core_sed_gates_record20_seqn;
assign main_genericstandalone_rtio_core_sed_record4_replace_occured = main_genericstandalone_rtio_core_sed_gates_record20_replace_occured;
assign main_genericstandalone_rtio_core_sed_record4_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record20_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record4_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record20_payload_channel;
assign main_genericstandalone_rtio_core_sed_record4_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record20_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record4_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record20_payload_address;
assign main_genericstandalone_rtio_core_sed_record4_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record20_payload_data;
assign main_genericstandalone_rtio_core_sed_record5_valid0 = main_genericstandalone_rtio_core_sed_gates_record21_valid;
assign main_genericstandalone_rtio_core_sed_record5_seqn1 = main_genericstandalone_rtio_core_sed_gates_record21_seqn;
assign main_genericstandalone_rtio_core_sed_record5_replace_occured = main_genericstandalone_rtio_core_sed_gates_record21_replace_occured;
assign main_genericstandalone_rtio_core_sed_record5_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record21_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record5_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record21_payload_channel;
assign main_genericstandalone_rtio_core_sed_record5_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record21_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record5_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record21_payload_address;
assign main_genericstandalone_rtio_core_sed_record5_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record21_payload_data;
assign main_genericstandalone_rtio_core_sed_record6_valid0 = main_genericstandalone_rtio_core_sed_gates_record22_valid;
assign main_genericstandalone_rtio_core_sed_record6_seqn1 = main_genericstandalone_rtio_core_sed_gates_record22_seqn;
assign main_genericstandalone_rtio_core_sed_record6_replace_occured = main_genericstandalone_rtio_core_sed_gates_record22_replace_occured;
assign main_genericstandalone_rtio_core_sed_record6_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record22_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record6_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record22_payload_channel;
assign main_genericstandalone_rtio_core_sed_record6_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record22_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record6_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record22_payload_address;
assign main_genericstandalone_rtio_core_sed_record6_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record22_payload_data;
assign main_genericstandalone_rtio_core_sed_record7_valid0 = main_genericstandalone_rtio_core_sed_gates_record23_valid;
assign main_genericstandalone_rtio_core_sed_record7_seqn1 = main_genericstandalone_rtio_core_sed_gates_record23_seqn;
assign main_genericstandalone_rtio_core_sed_record7_replace_occured = main_genericstandalone_rtio_core_sed_gates_record23_replace_occured;
assign main_genericstandalone_rtio_core_sed_record7_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record23_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record7_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record23_payload_channel;
assign main_genericstandalone_rtio_core_sed_record7_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record23_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record7_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record23_payload_address;
assign main_genericstandalone_rtio_core_sed_record7_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record23_payload_data;
assign main_genericstandalone_rtio_core_sed_record8_valid0 = main_genericstandalone_rtio_core_sed_gates_record24_valid;
assign main_genericstandalone_rtio_core_sed_record8_seqn1 = main_genericstandalone_rtio_core_sed_gates_record24_seqn;
assign main_genericstandalone_rtio_core_sed_record8_replace_occured = main_genericstandalone_rtio_core_sed_gates_record24_replace_occured;
assign main_genericstandalone_rtio_core_sed_record8_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record24_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record8_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record24_payload_channel;
assign main_genericstandalone_rtio_core_sed_record8_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record24_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record8_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record24_payload_address;
assign main_genericstandalone_rtio_core_sed_record8_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record24_payload_data;
assign main_genericstandalone_rtio_core_sed_record9_valid0 = main_genericstandalone_rtio_core_sed_gates_record25_valid;
assign main_genericstandalone_rtio_core_sed_record9_seqn1 = main_genericstandalone_rtio_core_sed_gates_record25_seqn;
assign main_genericstandalone_rtio_core_sed_record9_replace_occured = main_genericstandalone_rtio_core_sed_gates_record25_replace_occured;
assign main_genericstandalone_rtio_core_sed_record9_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record25_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record9_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record25_payload_channel;
assign main_genericstandalone_rtio_core_sed_record9_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record25_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record9_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record25_payload_address;
assign main_genericstandalone_rtio_core_sed_record9_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record25_payload_data;
assign main_genericstandalone_rtio_core_sed_record10_valid0 = main_genericstandalone_rtio_core_sed_gates_record26_valid;
assign main_genericstandalone_rtio_core_sed_record10_seqn1 = main_genericstandalone_rtio_core_sed_gates_record26_seqn;
assign main_genericstandalone_rtio_core_sed_record10_replace_occured = main_genericstandalone_rtio_core_sed_gates_record26_replace_occured;
assign main_genericstandalone_rtio_core_sed_record10_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record26_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record10_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record26_payload_channel;
assign main_genericstandalone_rtio_core_sed_record10_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record26_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record10_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record26_payload_address;
assign main_genericstandalone_rtio_core_sed_record10_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record26_payload_data;
assign main_genericstandalone_rtio_core_sed_record11_valid0 = main_genericstandalone_rtio_core_sed_gates_record27_valid;
assign main_genericstandalone_rtio_core_sed_record11_seqn1 = main_genericstandalone_rtio_core_sed_gates_record27_seqn;
assign main_genericstandalone_rtio_core_sed_record11_replace_occured = main_genericstandalone_rtio_core_sed_gates_record27_replace_occured;
assign main_genericstandalone_rtio_core_sed_record11_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record27_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record11_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record27_payload_channel;
assign main_genericstandalone_rtio_core_sed_record11_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record27_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record11_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record27_payload_address;
assign main_genericstandalone_rtio_core_sed_record11_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record27_payload_data;
assign main_genericstandalone_rtio_core_sed_record12_valid0 = main_genericstandalone_rtio_core_sed_gates_record28_valid;
assign main_genericstandalone_rtio_core_sed_record12_seqn1 = main_genericstandalone_rtio_core_sed_gates_record28_seqn;
assign main_genericstandalone_rtio_core_sed_record12_replace_occured = main_genericstandalone_rtio_core_sed_gates_record28_replace_occured;
assign main_genericstandalone_rtio_core_sed_record12_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record28_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record12_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record28_payload_channel;
assign main_genericstandalone_rtio_core_sed_record12_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record28_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record12_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record28_payload_address;
assign main_genericstandalone_rtio_core_sed_record12_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record28_payload_data;
assign main_genericstandalone_rtio_core_sed_record13_valid0 = main_genericstandalone_rtio_core_sed_gates_record29_valid;
assign main_genericstandalone_rtio_core_sed_record13_seqn1 = main_genericstandalone_rtio_core_sed_gates_record29_seqn;
assign main_genericstandalone_rtio_core_sed_record13_replace_occured = main_genericstandalone_rtio_core_sed_gates_record29_replace_occured;
assign main_genericstandalone_rtio_core_sed_record13_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record29_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record13_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record29_payload_channel;
assign main_genericstandalone_rtio_core_sed_record13_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record29_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record13_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record29_payload_address;
assign main_genericstandalone_rtio_core_sed_record13_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record29_payload_data;
assign main_genericstandalone_rtio_core_sed_record14_valid0 = main_genericstandalone_rtio_core_sed_gates_record30_valid;
assign main_genericstandalone_rtio_core_sed_record14_seqn1 = main_genericstandalone_rtio_core_sed_gates_record30_seqn;
assign main_genericstandalone_rtio_core_sed_record14_replace_occured = main_genericstandalone_rtio_core_sed_gates_record30_replace_occured;
assign main_genericstandalone_rtio_core_sed_record14_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record30_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record14_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record30_payload_channel;
assign main_genericstandalone_rtio_core_sed_record14_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record30_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record14_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record30_payload_address;
assign main_genericstandalone_rtio_core_sed_record14_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record30_payload_data;
assign main_genericstandalone_rtio_core_sed_record15_valid0 = main_genericstandalone_rtio_core_sed_gates_record31_valid;
assign main_genericstandalone_rtio_core_sed_record15_seqn1 = main_genericstandalone_rtio_core_sed_gates_record31_seqn;
assign main_genericstandalone_rtio_core_sed_record15_replace_occured = main_genericstandalone_rtio_core_sed_gates_record31_replace_occured;
assign main_genericstandalone_rtio_core_sed_record15_nondata_replace_occured = main_genericstandalone_rtio_core_sed_gates_record31_nondata_replace_occured;
assign main_genericstandalone_rtio_core_sed_record15_payload_channel1 = main_genericstandalone_rtio_core_sed_gates_record31_payload_channel;
assign main_genericstandalone_rtio_core_sed_record15_payload_fine_ts0 = main_genericstandalone_rtio_core_sed_gates_record31_payload_fine_ts;
assign main_genericstandalone_rtio_core_sed_record15_payload_address1 = main_genericstandalone_rtio_core_sed_gates_record31_payload_address;
assign main_genericstandalone_rtio_core_sed_record15_payload_data1 = main_genericstandalone_rtio_core_sed_gates_record31_payload_data;
assign main_genericstandalone_rtio_core_cri_o_status = {main_genericstandalone_rtio_core_sed_lane_dist_o_status_underflow, main_genericstandalone_rtio_core_sed_lane_dist_o_status_wait};
assign main_genericstandalone_rtio_core_sed_lane_dist_record0_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record1_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record2_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record3_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record4_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record5_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record6_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record7_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record8_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record9_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record10_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record11_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record12_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record13_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record14_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_record15_seqn = main_genericstandalone_rtio_core_sed_lane_dist_seqn;
assign main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_channel = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_address = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_data = main_genericstandalone_rtio_core_cri_o_data;
assign main_genericstandalone_rtio_core_sed_lane_dist_coarse_timestamp = main_genericstandalone_rtio_core_cri_o_timestamp[63:3];
assign main_genericstandalone_rtio_core_sed_lane_dist_current_lane_plus_one = (main_genericstandalone_rtio_core_sed_lane_dist_current_lane + 1'd1);
assign main_genericstandalone_rtio_core_sed_lane_dist_adr = main_genericstandalone_rtio_core_cri_chan_sel[15:0];
assign main_genericstandalone_rtio_core_sed_lane_dist_compensation = main_genericstandalone_rtio_core_sed_lane_dist_dat_r;
assign main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_min = ((main_genericstandalone_rtio_core_sed_lane_dist_min_minus_timestamp - main_genericstandalone_rtio_core_sed_lane_dist_compensation) < $signed({1'd0, 1'd0}));
assign main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_laneA_min = ((main_genericstandalone_rtio_core_sed_lane_dist_laneAmin_minus_timestamp - main_genericstandalone_rtio_core_sed_lane_dist_compensation) < $signed({1'd0, 1'd0}));
assign main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_laneB_min = ((main_genericstandalone_rtio_core_sed_lane_dist_laneBmin_minus_timestamp - main_genericstandalone_rtio_core_sed_lane_dist_compensation) < $signed({1'd0, 1'd0}));
assign main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_last = ((main_genericstandalone_rtio_core_sed_lane_dist_last_minus_timestamp - main_genericstandalone_rtio_core_sed_lane_dist_compensation) < $signed({1'd0, 1'd0}));

// synthesis translate_off
reg dummy_d_94;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_use_laneB <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_use_lanen <= 4'd0;
	if ((main_genericstandalone_rtio_core_sed_lane_dist_force_laneB | (~main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_last))) begin
		main_genericstandalone_rtio_core_sed_lane_dist_use_lanen <= main_genericstandalone_rtio_core_sed_lane_dist_current_lane_plus_one;
		main_genericstandalone_rtio_core_sed_lane_dist_use_laneB <= 1'd1;
	end else begin
		main_genericstandalone_rtio_core_sed_lane_dist_use_lanen <= main_genericstandalone_rtio_core_sed_lane_dist_current_lane;
		main_genericstandalone_rtio_core_sed_lane_dist_use_laneB <= 1'd0;
	end
// synthesis translate_off
	dummy_d_94 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_lane_min = (main_genericstandalone_rtio_core_sed_lane_dist_use_laneB ? main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_laneB_min : main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_laneA_min);

// synthesis translate_off
reg dummy_d_95;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_do_write <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_do_underflow <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_do_sequence_error <= 1'd0;
	if (((~main_genericstandalone_rtio_core_sed_lane_dist_quash) & (main_genericstandalone_rtio_core_cri_cmd == 1'd1))) begin
		if (main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_min) begin
			if (main_genericstandalone_rtio_core_sed_lane_dist_timestamp_above_lane_min) begin
				main_genericstandalone_rtio_core_sed_lane_dist_do_write <= 1'd1;
			end else begin
				main_genericstandalone_rtio_core_sed_lane_dist_do_sequence_error <= 1'd1;
			end
		end else begin
			main_genericstandalone_rtio_core_sed_lane_dist_do_underflow <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_95 <= dummy_s;
// synthesis translate_on
end
assign builder_comb_lhs_self = main_genericstandalone_rtio_core_sed_lane_dist_do_write;

// synthesis translate_off
reg dummy_d_96;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record0_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record1_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record2_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record3_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record4_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record5_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record6_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record7_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record8_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record9_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record10_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record11_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record12_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record13_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record14_we <= 1'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record15_we <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_lane_dist_use_lanen)
		1'd0: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record0_we <= builder_comb_lhs_self;
		end
		1'd1: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record1_we <= builder_comb_lhs_self;
		end
		2'd2: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record2_we <= builder_comb_lhs_self;
		end
		2'd3: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record3_we <= builder_comb_lhs_self;
		end
		3'd4: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record4_we <= builder_comb_lhs_self;
		end
		3'd5: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record5_we <= builder_comb_lhs_self;
		end
		3'd6: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record6_we <= builder_comb_lhs_self;
		end
		3'd7: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record7_we <= builder_comb_lhs_self;
		end
		4'd8: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record8_we <= builder_comb_lhs_self;
		end
		4'd9: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record9_we <= builder_comb_lhs_self;
		end
		4'd10: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record10_we <= builder_comb_lhs_self;
		end
		4'd11: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record11_we <= builder_comb_lhs_self;
		end
		4'd12: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record12_we <= builder_comb_lhs_self;
		end
		4'd13: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record13_we <= builder_comb_lhs_self;
		end
		4'd14: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record14_we <= builder_comb_lhs_self;
		end
		default: begin
			main_genericstandalone_rtio_core_sed_lane_dist_record15_we <= builder_comb_lhs_self;
		end
	endcase
// synthesis translate_off
	dummy_d_96 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp = ($signed({1'd0, main_genericstandalone_rtio_core_cri_o_timestamp}) + (main_genericstandalone_rtio_core_sed_lane_dist_compensation <<< 2'd3));

// synthesis translate_off
reg dummy_d_97;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record0_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_97 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_98;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record1_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_98 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_99;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record2_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_99 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_100;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record3_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_100 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_101;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record4_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_101 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_102;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record5_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_102 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_103;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record6_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_103 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_104;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record7_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_104 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_105;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record8_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_105 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_106;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record9_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_106 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_107;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record10_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_107 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_108;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record11_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_108 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_109;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record12_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_109 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_110;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record13_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_110 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_111;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record14_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_111 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_112;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_timestamp <= 64'd0;
	main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
	main_genericstandalone_rtio_core_sed_lane_dist_record15_payload_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp;
// synthesis translate_off
	dummy_d_112 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_lane_dist_current_lane_high_watermark = builder_comb_rhs_self8;
assign main_genericstandalone_rtio_core_sed_lane_dist_current_lane_writable = builder_comb_rhs_self9;
assign main_genericstandalone_rtio_core_sed_lane_dist_o_status_wait = (~main_genericstandalone_rtio_core_sed_lane_dist_current_lane_writable);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_din = {{main_genericstandalone_rtio_core_sed_record0_payload_data0, main_genericstandalone_rtio_core_sed_record0_payload_address0, main_genericstandalone_rtio_core_sed_record0_payload_timestamp, main_genericstandalone_rtio_core_sed_record0_payload_channel0}, main_genericstandalone_rtio_core_sed_record0_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_we = main_genericstandalone_rtio_core_sed_record0_we;
assign main_genericstandalone_rtio_core_sed_record0_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_writable;
assign main_genericstandalone_rtio_core_sed_record0_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered0_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record16_payload_data, main_genericstandalone_rtio_core_sed_record16_payload_address, main_genericstandalone_rtio_core_sed_record16_payload_timestamp, main_genericstandalone_rtio_core_sed_record16_payload_channel}, main_genericstandalone_rtio_core_sed_record16_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_dout;
assign main_genericstandalone_rtio_core_sed_record16_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered0_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_re = main_genericstandalone_rtio_core_sed_record16_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_din = {{main_genericstandalone_rtio_core_sed_record1_payload_data0, main_genericstandalone_rtio_core_sed_record1_payload_address0, main_genericstandalone_rtio_core_sed_record1_payload_timestamp, main_genericstandalone_rtio_core_sed_record1_payload_channel0}, main_genericstandalone_rtio_core_sed_record1_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_we = main_genericstandalone_rtio_core_sed_record1_we;
assign main_genericstandalone_rtio_core_sed_record1_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_writable;
assign main_genericstandalone_rtio_core_sed_record1_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered1_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record17_payload_data, main_genericstandalone_rtio_core_sed_record17_payload_address, main_genericstandalone_rtio_core_sed_record17_payload_timestamp, main_genericstandalone_rtio_core_sed_record17_payload_channel}, main_genericstandalone_rtio_core_sed_record17_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_dout;
assign main_genericstandalone_rtio_core_sed_record17_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered1_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_re = main_genericstandalone_rtio_core_sed_record17_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_din = {{main_genericstandalone_rtio_core_sed_record2_payload_data0, main_genericstandalone_rtio_core_sed_record2_payload_address0, main_genericstandalone_rtio_core_sed_record2_payload_timestamp, main_genericstandalone_rtio_core_sed_record2_payload_channel0}, main_genericstandalone_rtio_core_sed_record2_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_we = main_genericstandalone_rtio_core_sed_record2_we;
assign main_genericstandalone_rtio_core_sed_record2_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_writable;
assign main_genericstandalone_rtio_core_sed_record2_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered2_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record18_payload_data, main_genericstandalone_rtio_core_sed_record18_payload_address, main_genericstandalone_rtio_core_sed_record18_payload_timestamp, main_genericstandalone_rtio_core_sed_record18_payload_channel}, main_genericstandalone_rtio_core_sed_record18_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_dout;
assign main_genericstandalone_rtio_core_sed_record18_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered2_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_re = main_genericstandalone_rtio_core_sed_record18_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_din = {{main_genericstandalone_rtio_core_sed_record3_payload_data0, main_genericstandalone_rtio_core_sed_record3_payload_address0, main_genericstandalone_rtio_core_sed_record3_payload_timestamp, main_genericstandalone_rtio_core_sed_record3_payload_channel0}, main_genericstandalone_rtio_core_sed_record3_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_we = main_genericstandalone_rtio_core_sed_record3_we;
assign main_genericstandalone_rtio_core_sed_record3_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_writable;
assign main_genericstandalone_rtio_core_sed_record3_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered3_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record19_payload_data, main_genericstandalone_rtio_core_sed_record19_payload_address, main_genericstandalone_rtio_core_sed_record19_payload_timestamp, main_genericstandalone_rtio_core_sed_record19_payload_channel}, main_genericstandalone_rtio_core_sed_record19_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_dout;
assign main_genericstandalone_rtio_core_sed_record19_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered3_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_re = main_genericstandalone_rtio_core_sed_record19_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_din = {{main_genericstandalone_rtio_core_sed_record4_payload_data0, main_genericstandalone_rtio_core_sed_record4_payload_address0, main_genericstandalone_rtio_core_sed_record4_payload_timestamp, main_genericstandalone_rtio_core_sed_record4_payload_channel0}, main_genericstandalone_rtio_core_sed_record4_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_we = main_genericstandalone_rtio_core_sed_record4_we;
assign main_genericstandalone_rtio_core_sed_record4_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_writable;
assign main_genericstandalone_rtio_core_sed_record4_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered4_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record20_payload_data, main_genericstandalone_rtio_core_sed_record20_payload_address, main_genericstandalone_rtio_core_sed_record20_payload_timestamp, main_genericstandalone_rtio_core_sed_record20_payload_channel}, main_genericstandalone_rtio_core_sed_record20_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_dout;
assign main_genericstandalone_rtio_core_sed_record20_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered4_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_re = main_genericstandalone_rtio_core_sed_record20_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_din = {{main_genericstandalone_rtio_core_sed_record5_payload_data0, main_genericstandalone_rtio_core_sed_record5_payload_address0, main_genericstandalone_rtio_core_sed_record5_payload_timestamp, main_genericstandalone_rtio_core_sed_record5_payload_channel0}, main_genericstandalone_rtio_core_sed_record5_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_we = main_genericstandalone_rtio_core_sed_record5_we;
assign main_genericstandalone_rtio_core_sed_record5_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_writable;
assign main_genericstandalone_rtio_core_sed_record5_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered5_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record21_payload_data, main_genericstandalone_rtio_core_sed_record21_payload_address, main_genericstandalone_rtio_core_sed_record21_payload_timestamp, main_genericstandalone_rtio_core_sed_record21_payload_channel}, main_genericstandalone_rtio_core_sed_record21_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_dout;
assign main_genericstandalone_rtio_core_sed_record21_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered5_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_re = main_genericstandalone_rtio_core_sed_record21_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_din = {{main_genericstandalone_rtio_core_sed_record6_payload_data0, main_genericstandalone_rtio_core_sed_record6_payload_address0, main_genericstandalone_rtio_core_sed_record6_payload_timestamp, main_genericstandalone_rtio_core_sed_record6_payload_channel0}, main_genericstandalone_rtio_core_sed_record6_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_we = main_genericstandalone_rtio_core_sed_record6_we;
assign main_genericstandalone_rtio_core_sed_record6_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_writable;
assign main_genericstandalone_rtio_core_sed_record6_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered6_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record22_payload_data, main_genericstandalone_rtio_core_sed_record22_payload_address, main_genericstandalone_rtio_core_sed_record22_payload_timestamp, main_genericstandalone_rtio_core_sed_record22_payload_channel}, main_genericstandalone_rtio_core_sed_record22_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_dout;
assign main_genericstandalone_rtio_core_sed_record22_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered6_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_re = main_genericstandalone_rtio_core_sed_record22_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_din = {{main_genericstandalone_rtio_core_sed_record7_payload_data0, main_genericstandalone_rtio_core_sed_record7_payload_address0, main_genericstandalone_rtio_core_sed_record7_payload_timestamp, main_genericstandalone_rtio_core_sed_record7_payload_channel0}, main_genericstandalone_rtio_core_sed_record7_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_we = main_genericstandalone_rtio_core_sed_record7_we;
assign main_genericstandalone_rtio_core_sed_record7_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_writable;
assign main_genericstandalone_rtio_core_sed_record7_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered7_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record23_payload_data, main_genericstandalone_rtio_core_sed_record23_payload_address, main_genericstandalone_rtio_core_sed_record23_payload_timestamp, main_genericstandalone_rtio_core_sed_record23_payload_channel}, main_genericstandalone_rtio_core_sed_record23_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_dout;
assign main_genericstandalone_rtio_core_sed_record23_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered7_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_re = main_genericstandalone_rtio_core_sed_record23_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_din = {{main_genericstandalone_rtio_core_sed_record8_payload_data0, main_genericstandalone_rtio_core_sed_record8_payload_address0, main_genericstandalone_rtio_core_sed_record8_payload_timestamp, main_genericstandalone_rtio_core_sed_record8_payload_channel0}, main_genericstandalone_rtio_core_sed_record8_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_we = main_genericstandalone_rtio_core_sed_record8_we;
assign main_genericstandalone_rtio_core_sed_record8_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_writable;
assign main_genericstandalone_rtio_core_sed_record8_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered8_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record24_payload_data, main_genericstandalone_rtio_core_sed_record24_payload_address, main_genericstandalone_rtio_core_sed_record24_payload_timestamp, main_genericstandalone_rtio_core_sed_record24_payload_channel}, main_genericstandalone_rtio_core_sed_record24_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_dout;
assign main_genericstandalone_rtio_core_sed_record24_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered8_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_re = main_genericstandalone_rtio_core_sed_record24_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_din = {{main_genericstandalone_rtio_core_sed_record9_payload_data0, main_genericstandalone_rtio_core_sed_record9_payload_address0, main_genericstandalone_rtio_core_sed_record9_payload_timestamp, main_genericstandalone_rtio_core_sed_record9_payload_channel0}, main_genericstandalone_rtio_core_sed_record9_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_we = main_genericstandalone_rtio_core_sed_record9_we;
assign main_genericstandalone_rtio_core_sed_record9_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_writable;
assign main_genericstandalone_rtio_core_sed_record9_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered9_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record25_payload_data, main_genericstandalone_rtio_core_sed_record25_payload_address, main_genericstandalone_rtio_core_sed_record25_payload_timestamp, main_genericstandalone_rtio_core_sed_record25_payload_channel}, main_genericstandalone_rtio_core_sed_record25_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_dout;
assign main_genericstandalone_rtio_core_sed_record25_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered9_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_re = main_genericstandalone_rtio_core_sed_record25_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_din = {{main_genericstandalone_rtio_core_sed_record10_payload_data0, main_genericstandalone_rtio_core_sed_record10_payload_address0, main_genericstandalone_rtio_core_sed_record10_payload_timestamp, main_genericstandalone_rtio_core_sed_record10_payload_channel0}, main_genericstandalone_rtio_core_sed_record10_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_we = main_genericstandalone_rtio_core_sed_record10_we;
assign main_genericstandalone_rtio_core_sed_record10_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_writable;
assign main_genericstandalone_rtio_core_sed_record10_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered10_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record26_payload_data, main_genericstandalone_rtio_core_sed_record26_payload_address, main_genericstandalone_rtio_core_sed_record26_payload_timestamp, main_genericstandalone_rtio_core_sed_record26_payload_channel}, main_genericstandalone_rtio_core_sed_record26_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_dout;
assign main_genericstandalone_rtio_core_sed_record26_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered10_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_re = main_genericstandalone_rtio_core_sed_record26_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_din = {{main_genericstandalone_rtio_core_sed_record11_payload_data0, main_genericstandalone_rtio_core_sed_record11_payload_address0, main_genericstandalone_rtio_core_sed_record11_payload_timestamp, main_genericstandalone_rtio_core_sed_record11_payload_channel0}, main_genericstandalone_rtio_core_sed_record11_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_we = main_genericstandalone_rtio_core_sed_record11_we;
assign main_genericstandalone_rtio_core_sed_record11_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_writable;
assign main_genericstandalone_rtio_core_sed_record11_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered11_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record27_payload_data, main_genericstandalone_rtio_core_sed_record27_payload_address, main_genericstandalone_rtio_core_sed_record27_payload_timestamp, main_genericstandalone_rtio_core_sed_record27_payload_channel}, main_genericstandalone_rtio_core_sed_record27_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_dout;
assign main_genericstandalone_rtio_core_sed_record27_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered11_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_re = main_genericstandalone_rtio_core_sed_record27_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_din = {{main_genericstandalone_rtio_core_sed_record12_payload_data0, main_genericstandalone_rtio_core_sed_record12_payload_address0, main_genericstandalone_rtio_core_sed_record12_payload_timestamp, main_genericstandalone_rtio_core_sed_record12_payload_channel0}, main_genericstandalone_rtio_core_sed_record12_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_we = main_genericstandalone_rtio_core_sed_record12_we;
assign main_genericstandalone_rtio_core_sed_record12_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_writable;
assign main_genericstandalone_rtio_core_sed_record12_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered12_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record28_payload_data, main_genericstandalone_rtio_core_sed_record28_payload_address, main_genericstandalone_rtio_core_sed_record28_payload_timestamp, main_genericstandalone_rtio_core_sed_record28_payload_channel}, main_genericstandalone_rtio_core_sed_record28_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_dout;
assign main_genericstandalone_rtio_core_sed_record28_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered12_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_re = main_genericstandalone_rtio_core_sed_record28_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_din = {{main_genericstandalone_rtio_core_sed_record13_payload_data0, main_genericstandalone_rtio_core_sed_record13_payload_address0, main_genericstandalone_rtio_core_sed_record13_payload_timestamp, main_genericstandalone_rtio_core_sed_record13_payload_channel0}, main_genericstandalone_rtio_core_sed_record13_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_we = main_genericstandalone_rtio_core_sed_record13_we;
assign main_genericstandalone_rtio_core_sed_record13_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_writable;
assign main_genericstandalone_rtio_core_sed_record13_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered13_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record29_payload_data, main_genericstandalone_rtio_core_sed_record29_payload_address, main_genericstandalone_rtio_core_sed_record29_payload_timestamp, main_genericstandalone_rtio_core_sed_record29_payload_channel}, main_genericstandalone_rtio_core_sed_record29_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_dout;
assign main_genericstandalone_rtio_core_sed_record29_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered13_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_re = main_genericstandalone_rtio_core_sed_record29_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_din = {{main_genericstandalone_rtio_core_sed_record14_payload_data0, main_genericstandalone_rtio_core_sed_record14_payload_address0, main_genericstandalone_rtio_core_sed_record14_payload_timestamp, main_genericstandalone_rtio_core_sed_record14_payload_channel0}, main_genericstandalone_rtio_core_sed_record14_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_we = main_genericstandalone_rtio_core_sed_record14_we;
assign main_genericstandalone_rtio_core_sed_record14_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_writable;
assign main_genericstandalone_rtio_core_sed_record14_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered14_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record30_payload_data, main_genericstandalone_rtio_core_sed_record30_payload_address, main_genericstandalone_rtio_core_sed_record30_payload_timestamp, main_genericstandalone_rtio_core_sed_record30_payload_channel}, main_genericstandalone_rtio_core_sed_record30_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_dout;
assign main_genericstandalone_rtio_core_sed_record30_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered14_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_re = main_genericstandalone_rtio_core_sed_record30_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_din = {{main_genericstandalone_rtio_core_sed_record15_payload_data0, main_genericstandalone_rtio_core_sed_record15_payload_address0, main_genericstandalone_rtio_core_sed_record15_payload_timestamp, main_genericstandalone_rtio_core_sed_record15_payload_channel0}, main_genericstandalone_rtio_core_sed_record15_seqn0};
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_we = main_genericstandalone_rtio_core_sed_record15_we;
assign main_genericstandalone_rtio_core_sed_record15_writable = main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_writable;
assign main_genericstandalone_rtio_core_sed_record15_high_watermark = (main_genericstandalone_rtio_core_sed_syncfifobuffered15_level1 >= 8'd128);
assign {{main_genericstandalone_rtio_core_sed_record31_payload_data, main_genericstandalone_rtio_core_sed_record31_payload_address, main_genericstandalone_rtio_core_sed_record31_payload_timestamp, main_genericstandalone_rtio_core_sed_record31_payload_channel}, main_genericstandalone_rtio_core_sed_record31_seqn} = main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_dout;
assign main_genericstandalone_rtio_core_sed_record31_readable = main_genericstandalone_rtio_core_sed_syncfifobuffered15_readable;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_re = main_genericstandalone_rtio_core_sed_record31_re;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered0_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered0_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered0_readable);

// synthesis translate_off
reg dummy_d_113;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered0_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered0_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered0_produce;
	end
// synthesis translate_off
	dummy_d_113 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered0_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered0_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered0_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered1_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered1_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered1_readable);

// synthesis translate_off
reg dummy_d_114;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered1_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered1_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered1_produce;
	end
// synthesis translate_off
	dummy_d_114 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered1_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered1_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered1_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered2_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered2_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered2_readable);

// synthesis translate_off
reg dummy_d_115;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered2_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered2_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered2_produce;
	end
// synthesis translate_off
	dummy_d_115 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered2_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered2_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered2_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered3_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered3_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered3_readable);

// synthesis translate_off
reg dummy_d_116;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered3_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered3_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered3_produce;
	end
// synthesis translate_off
	dummy_d_116 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered3_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered3_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered3_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered4_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered4_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered4_readable);

// synthesis translate_off
reg dummy_d_117;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered4_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered4_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered4_produce;
	end
// synthesis translate_off
	dummy_d_117 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered4_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered4_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered4_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered5_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered5_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered5_readable);

// synthesis translate_off
reg dummy_d_118;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered5_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered5_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered5_produce;
	end
// synthesis translate_off
	dummy_d_118 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered5_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered5_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered5_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered6_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered6_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered6_readable);

// synthesis translate_off
reg dummy_d_119;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered6_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered6_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered6_produce;
	end
// synthesis translate_off
	dummy_d_119 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered6_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered6_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered6_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered7_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered7_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered7_readable);

// synthesis translate_off
reg dummy_d_120;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered7_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered7_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered7_produce;
	end
// synthesis translate_off
	dummy_d_120 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered7_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered7_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered7_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered8_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered8_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered8_readable);

// synthesis translate_off
reg dummy_d_121;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered8_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered8_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered8_produce;
	end
// synthesis translate_off
	dummy_d_121 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered8_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered8_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered8_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered9_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered9_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered9_readable);

// synthesis translate_off
reg dummy_d_122;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered9_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered9_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered9_produce;
	end
// synthesis translate_off
	dummy_d_122 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered9_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered9_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered9_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered10_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered10_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered10_readable);

// synthesis translate_off
reg dummy_d_123;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered10_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered10_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered10_produce;
	end
// synthesis translate_off
	dummy_d_123 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered10_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered10_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered10_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered11_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered11_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered11_readable);

// synthesis translate_off
reg dummy_d_124;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered11_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered11_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered11_produce;
	end
// synthesis translate_off
	dummy_d_124 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered11_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered11_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered11_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered12_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered12_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered12_readable);

// synthesis translate_off
reg dummy_d_125;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered12_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered12_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered12_produce;
	end
// synthesis translate_off
	dummy_d_125 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered12_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered12_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered12_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered13_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered13_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered13_readable);

// synthesis translate_off
reg dummy_d_126;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered13_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered13_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered13_produce;
	end
// synthesis translate_off
	dummy_d_126 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered13_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered13_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered13_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered14_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered14_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered14_readable);

// synthesis translate_off
reg dummy_d_127;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered14_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered14_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered14_produce;
	end
// synthesis translate_off
	dummy_d_127 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered14_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered14_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered14_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_re = (main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_readable & ((~main_genericstandalone_rtio_core_sed_syncfifobuffered15_readable) | main_genericstandalone_rtio_core_sed_syncfifobuffered15_re));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_level1 = (main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 + main_genericstandalone_rtio_core_sed_syncfifobuffered15_readable);

// synthesis translate_off
reg dummy_d_128;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered15_replace) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_adr <= (main_genericstandalone_rtio_core_sed_syncfifobuffered15_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_adr <= main_genericstandalone_rtio_core_sed_syncfifobuffered15_produce;
	end
// synthesis translate_off
	dummy_d_128 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_dat_w = main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_din;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_we = (main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_we & (main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_writable | main_genericstandalone_rtio_core_sed_syncfifobuffered15_replace));
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_do_read = (main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_readable & main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_re);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_adr = main_genericstandalone_rtio_core_sed_syncfifobuffered15_consume;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_dout = main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_dat_r;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_re = main_genericstandalone_rtio_core_sed_syncfifobuffered15_do_read;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_writable = (main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 != 8'd128);
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_readable = (main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 != 1'd0);
assign main_genericstandalone_rtio_core_sed_gates_record16_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record16_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record0_re = (main_genericstandalone_rtio_core_sed_gates_record0_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record17_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record17_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record1_re = (main_genericstandalone_rtio_core_sed_gates_record1_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record18_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record18_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record2_re = (main_genericstandalone_rtio_core_sed_gates_record2_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record19_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record19_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record3_re = (main_genericstandalone_rtio_core_sed_gates_record3_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record20_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record20_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record4_re = (main_genericstandalone_rtio_core_sed_gates_record4_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record21_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record21_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record5_re = (main_genericstandalone_rtio_core_sed_gates_record5_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record22_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record22_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record6_re = (main_genericstandalone_rtio_core_sed_gates_record6_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record23_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record23_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record7_re = (main_genericstandalone_rtio_core_sed_gates_record7_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record24_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record24_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record8_re = (main_genericstandalone_rtio_core_sed_gates_record8_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record25_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record25_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record9_re = (main_genericstandalone_rtio_core_sed_gates_record9_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record26_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record26_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record10_re = (main_genericstandalone_rtio_core_sed_gates_record10_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record27_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record27_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record11_re = (main_genericstandalone_rtio_core_sed_gates_record11_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record28_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record28_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record12_re = (main_genericstandalone_rtio_core_sed_gates_record12_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record29_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record29_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record13_re = (main_genericstandalone_rtio_core_sed_gates_record13_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record30_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record30_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record14_re = (main_genericstandalone_rtio_core_sed_gates_record14_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_gates_record31_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record31_nondata_replace_occured = 1'd0;
assign main_genericstandalone_rtio_core_sed_gates_record15_re = (main_genericstandalone_rtio_core_sed_gates_record15_payload_timestamp[63:3] == main_genericstandalone_rtio_core_sed_gates_coarse_timestamp);
assign main_genericstandalone_rtio_core_sed_memory0_adr = main_genericstandalone_rtio_core_sed_record144_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record0_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r0 & ((~main_genericstandalone_rtio_core_sed_memory0_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r0));
assign main_genericstandalone_rtio_core_sed_memory1_adr = main_genericstandalone_rtio_core_sed_record145_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record1_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r1 & ((~main_genericstandalone_rtio_core_sed_memory1_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r1));
assign main_genericstandalone_rtio_core_sed_memory2_adr = main_genericstandalone_rtio_core_sed_record146_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record2_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r2 & ((~main_genericstandalone_rtio_core_sed_memory2_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r2));
assign main_genericstandalone_rtio_core_sed_memory3_adr = main_genericstandalone_rtio_core_sed_record147_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record3_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r3 & ((~main_genericstandalone_rtio_core_sed_memory3_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r3));
assign main_genericstandalone_rtio_core_sed_memory4_adr = main_genericstandalone_rtio_core_sed_record148_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record4_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r4 & ((~main_genericstandalone_rtio_core_sed_memory4_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r4));
assign main_genericstandalone_rtio_core_sed_memory5_adr = main_genericstandalone_rtio_core_sed_record149_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record5_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r5 & ((~main_genericstandalone_rtio_core_sed_memory5_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r5));
assign main_genericstandalone_rtio_core_sed_memory6_adr = main_genericstandalone_rtio_core_sed_record150_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record6_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r6 & ((~main_genericstandalone_rtio_core_sed_memory6_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r6));
assign main_genericstandalone_rtio_core_sed_memory7_adr = main_genericstandalone_rtio_core_sed_record151_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record7_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r7 & ((~main_genericstandalone_rtio_core_sed_memory7_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r7));
assign main_genericstandalone_rtio_core_sed_memory8_adr = main_genericstandalone_rtio_core_sed_record152_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record8_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r8 & ((~main_genericstandalone_rtio_core_sed_memory8_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r8));
assign main_genericstandalone_rtio_core_sed_memory9_adr = main_genericstandalone_rtio_core_sed_record153_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record9_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r9 & ((~main_genericstandalone_rtio_core_sed_memory9_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r9));
assign main_genericstandalone_rtio_core_sed_memory10_adr = main_genericstandalone_rtio_core_sed_record154_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record10_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r10 & ((~main_genericstandalone_rtio_core_sed_memory10_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r10));
assign main_genericstandalone_rtio_core_sed_memory11_adr = main_genericstandalone_rtio_core_sed_record155_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record11_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r11 & ((~main_genericstandalone_rtio_core_sed_memory11_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r11));
assign main_genericstandalone_rtio_core_sed_memory12_adr = main_genericstandalone_rtio_core_sed_record156_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record12_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r12 & ((~main_genericstandalone_rtio_core_sed_memory12_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r12));
assign main_genericstandalone_rtio_core_sed_memory13_adr = main_genericstandalone_rtio_core_sed_record157_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record13_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r13 & ((~main_genericstandalone_rtio_core_sed_memory13_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r13));
assign main_genericstandalone_rtio_core_sed_memory14_adr = main_genericstandalone_rtio_core_sed_record158_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record14_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r14 & ((~main_genericstandalone_rtio_core_sed_memory14_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r14));
assign main_genericstandalone_rtio_core_sed_memory15_adr = main_genericstandalone_rtio_core_sed_record159_rec_payload_channel;
assign main_genericstandalone_rtio_core_sed_record15_collision = (main_genericstandalone_rtio_core_sed_replace_occured_r15 & ((~main_genericstandalone_rtio_core_sed_memory15_dat_r) | main_genericstandalone_rtio_core_sed_nondata_replace_occured_r15));
assign main_genericstandalone_rtio_core_sed_selected0 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected1 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected2 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected3 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected4 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected5 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected6 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected7 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected8 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected9 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected10 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected11 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected12 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected13 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected14 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected15 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 1'd0));
assign main_genericstandalone_rtio_core_sed_selected16 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected17 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected18 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected19 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected20 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected21 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected22 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected23 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected24 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected25 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected26 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected27 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected28 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected29 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected30 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected31 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 1'd1));
assign main_genericstandalone_rtio_core_sed_selected32 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected33 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected34 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected35 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected36 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected37 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected38 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected39 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected40 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected41 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected42 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected43 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected44 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected45 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected46 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected47 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 2'd2));
assign main_genericstandalone_rtio_core_sed_selected48 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected49 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected50 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected51 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected52 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected53 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected54 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected55 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected56 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected57 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected58 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected59 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected60 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected61 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected62 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected63 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 2'd3));
assign main_genericstandalone_rtio_core_sed_selected64 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected65 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected66 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected67 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected68 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected69 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected70 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected71 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected72 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected73 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected74 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected75 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected76 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected77 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected78 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected79 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 3'd4));
assign main_genericstandalone_rtio_core_sed_selected80 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected81 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected82 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected83 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected84 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected85 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected86 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected87 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected88 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected89 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected90 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected91 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected92 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected93 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected94 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected95 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 3'd5));
assign main_genericstandalone_rtio_core_sed_selected96 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected97 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected98 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected99 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected100 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected101 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected102 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected103 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected104 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected105 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected106 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected107 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected108 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected109 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected110 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected111 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 3'd6));
assign main_genericstandalone_rtio_core_sed_selected112 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected113 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected114 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected115 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected116 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected117 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected118 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected119 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected120 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected121 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected122 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected123 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected124 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected125 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected126 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected127 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 3'd7));
assign main_genericstandalone_rtio_core_sed_selected128 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected129 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected130 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected131 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected132 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected133 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected134 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected135 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected136 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected137 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected138 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected139 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected140 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected141 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected142 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected143 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 4'd8));
assign main_genericstandalone_rtio_core_sed_selected144 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected145 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected146 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected147 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected148 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected149 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected150 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected151 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected152 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected153 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected154 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected155 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected156 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected157 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected158 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected159 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 4'd9));
assign main_genericstandalone_rtio_core_sed_selected160 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected161 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected162 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected163 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected164 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected165 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected166 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected167 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected168 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected169 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected170 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected171 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected172 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected173 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected174 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected175 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 4'd10));
assign main_genericstandalone_rtio_core_sed_selected176 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected177 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected178 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected179 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected180 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected181 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected182 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected183 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected184 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected185 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected186 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected187 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected188 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected189 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected190 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected191 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 4'd11));
assign main_genericstandalone_rtio_core_sed_selected192 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected193 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected194 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected195 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected196 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected197 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected198 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected199 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected200 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected201 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected202 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected203 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected204 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected205 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected206 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected207 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 4'd12));
assign main_genericstandalone_rtio_core_sed_selected208 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected209 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected210 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected211 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected212 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected213 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected214 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected215 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected216 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected217 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected218 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected219 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected220 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected221 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected222 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected223 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 4'd13));
assign main_genericstandalone_rtio_core_sed_selected224 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected225 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected226 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected227 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected228 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected229 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected230 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected231 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected232 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected233 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected234 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected235 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected236 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected237 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected238 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected239 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 4'd14));
assign main_genericstandalone_rtio_core_sed_selected240 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected241 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected242 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected243 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected244 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected245 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected246 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected247 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected248 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected249 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected250 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected251 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected252 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected253 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected254 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected255 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 4'd15));
assign main_genericstandalone_rtio_core_sed_selected256 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected257 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected258 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected259 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected260 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected261 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected262 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected263 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected264 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected265 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected266 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected267 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected268 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected269 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected270 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected271 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd16));
assign main_genericstandalone_rtio_core_sed_selected272 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected273 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected274 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected275 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected276 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected277 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected278 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected279 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected280 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected281 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected282 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected283 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected284 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected285 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected286 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected287 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd17));
assign main_genericstandalone_rtio_core_sed_selected288 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected289 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected290 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected291 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected292 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected293 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected294 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected295 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected296 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected297 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected298 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected299 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected300 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected301 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected302 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected303 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd18));
assign main_genericstandalone_rtio_core_sed_selected304 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected305 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected306 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected307 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected308 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected309 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected310 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected311 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected312 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected313 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected314 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected315 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected316 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected317 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected318 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected319 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd19));
assign main_genericstandalone_rtio_core_sed_selected320 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected321 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected322 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected323 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected324 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected325 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected326 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected327 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected328 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected329 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected330 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected331 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected332 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected333 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected334 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected335 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd20));
assign main_genericstandalone_rtio_core_sed_selected336 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected337 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected338 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected339 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected340 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected341 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected342 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected343 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected344 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected345 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected346 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected347 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected348 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected349 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected350 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected351 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd21));
assign main_genericstandalone_rtio_core_sed_selected352 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected353 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected354 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected355 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected356 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected357 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected358 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected359 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected360 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected361 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected362 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected363 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected364 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected365 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected366 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected367 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd22));
assign main_genericstandalone_rtio_core_sed_selected368 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected369 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected370 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected371 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected372 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected373 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected374 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected375 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected376 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected377 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected378 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected379 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected380 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected381 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected382 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected383 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd23));
assign main_genericstandalone_rtio_core_sed_selected384 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected385 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected386 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected387 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected388 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected389 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected390 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected391 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected392 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected393 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected394 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected395 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected396 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected397 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected398 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected399 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd24));
assign main_genericstandalone_rtio_core_sed_selected400 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected401 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected402 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected403 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected404 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected405 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected406 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected407 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected408 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected409 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected410 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected411 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected412 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected413 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected414 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected415 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd25));
assign main_genericstandalone_rtio_core_sed_selected416 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected417 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected418 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected419 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected420 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected421 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected422 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected423 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected424 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected425 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected426 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected427 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected428 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected429 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected430 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected431 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd26));
assign main_genericstandalone_rtio_core_sed_selected432 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected433 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected434 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected435 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected436 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected437 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected438 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected439 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected440 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected441 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected442 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected443 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected444 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected445 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected446 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected447 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd27));
assign main_genericstandalone_rtio_core_sed_selected448 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected449 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected450 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected451 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected452 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected453 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected454 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected455 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected456 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected457 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected458 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected459 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected460 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected461 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected462 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected463 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd28));
assign main_genericstandalone_rtio_core_sed_selected464 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected465 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected466 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected467 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected468 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected469 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected470 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected471 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected472 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected473 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected474 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected475 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected476 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected477 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected478 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected479 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd29));
assign main_genericstandalone_rtio_core_sed_selected480 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected481 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected482 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected483 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected484 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected485 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected486 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected487 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected488 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected489 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected490 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected491 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected492 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected493 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected494 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected495 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd30));
assign main_genericstandalone_rtio_core_sed_selected496 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected497 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected498 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected499 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected500 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected501 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected502 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected503 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected504 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected505 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected506 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected507 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected508 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected509 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected510 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected511 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 5'd31));
assign main_genericstandalone_rtio_core_sed_selected512 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected513 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected514 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected515 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected516 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected517 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected518 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected519 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected520 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected521 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected522 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected523 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected524 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected525 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected526 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected527 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 6'd32));
assign main_genericstandalone_rtio_core_sed_selected528 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected529 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected530 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected531 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected532 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected533 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected534 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected535 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected536 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected537 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected538 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected539 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected540 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected541 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected542 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected543 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 6'd33));
assign main_genericstandalone_rtio_core_sed_selected544 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected545 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected546 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected547 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected548 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected549 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected550 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected551 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected552 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected553 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected554 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected555 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected556 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected557 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected558 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected559 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 6'd34));
assign main_genericstandalone_rtio_core_sed_selected560 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected561 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected562 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected563 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected564 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected565 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected566 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected567 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected568 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected569 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected570 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected571 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected572 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected573 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected574 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected575 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 6'd35));
assign main_genericstandalone_rtio_core_sed_selected576 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected577 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected578 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected579 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected580 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected581 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected582 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected583 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected584 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected585 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected586 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected587 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected588 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected589 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected590 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected591 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 6'd36));
assign main_genericstandalone_rtio_core_sed_selected592 = ((main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision)) & (main_genericstandalone_rtio_core_sed_record0_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected593 = ((main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision)) & (main_genericstandalone_rtio_core_sed_record1_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected594 = ((main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision)) & (main_genericstandalone_rtio_core_sed_record2_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected595 = ((main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision)) & (main_genericstandalone_rtio_core_sed_record3_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected596 = ((main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision)) & (main_genericstandalone_rtio_core_sed_record4_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected597 = ((main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision)) & (main_genericstandalone_rtio_core_sed_record5_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected598 = ((main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision)) & (main_genericstandalone_rtio_core_sed_record6_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected599 = ((main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision)) & (main_genericstandalone_rtio_core_sed_record7_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected600 = ((main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision)) & (main_genericstandalone_rtio_core_sed_record8_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected601 = ((main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision)) & (main_genericstandalone_rtio_core_sed_record9_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected602 = ((main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision)) & (main_genericstandalone_rtio_core_sed_record10_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected603 = ((main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision)) & (main_genericstandalone_rtio_core_sed_record11_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected604 = ((main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision)) & (main_genericstandalone_rtio_core_sed_record12_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected605 = ((main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision)) & (main_genericstandalone_rtio_core_sed_record13_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected606 = ((main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision)) & (main_genericstandalone_rtio_core_sed_record14_payload_channel2 == 6'd37));
assign main_genericstandalone_rtio_core_sed_selected607 = ((main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision)) & (main_genericstandalone_rtio_core_sed_record15_payload_channel2 == 6'd37));

// synthesis translate_off
reg dummy_d_129;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference0 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record0_payload_channel1 != main_genericstandalone_rtio_core_sed_record1_payload_channel1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference0 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record0_payload_fine_ts0 != main_genericstandalone_rtio_core_sed_record1_payload_fine_ts0)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference0 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record0_payload_address1 != main_genericstandalone_rtio_core_sed_record1_payload_address1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference0 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_129 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_130;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference1 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record2_payload_channel1 != main_genericstandalone_rtio_core_sed_record3_payload_channel1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference1 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record2_payload_fine_ts0 != main_genericstandalone_rtio_core_sed_record3_payload_fine_ts0)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference1 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record2_payload_address1 != main_genericstandalone_rtio_core_sed_record3_payload_address1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference1 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_130 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_131;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference2 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record4_payload_channel1 != main_genericstandalone_rtio_core_sed_record5_payload_channel1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference2 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record4_payload_fine_ts0 != main_genericstandalone_rtio_core_sed_record5_payload_fine_ts0)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference2 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record4_payload_address1 != main_genericstandalone_rtio_core_sed_record5_payload_address1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference2 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_131 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_132;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference3 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record6_payload_channel1 != main_genericstandalone_rtio_core_sed_record7_payload_channel1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference3 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record6_payload_fine_ts0 != main_genericstandalone_rtio_core_sed_record7_payload_fine_ts0)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference3 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record6_payload_address1 != main_genericstandalone_rtio_core_sed_record7_payload_address1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference3 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_132 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_133;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference4 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record8_payload_channel1 != main_genericstandalone_rtio_core_sed_record9_payload_channel1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference4 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record8_payload_fine_ts0 != main_genericstandalone_rtio_core_sed_record9_payload_fine_ts0)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference4 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record8_payload_address1 != main_genericstandalone_rtio_core_sed_record9_payload_address1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference4 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_133 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_134;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference5 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record10_payload_channel1 != main_genericstandalone_rtio_core_sed_record11_payload_channel1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference5 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record10_payload_fine_ts0 != main_genericstandalone_rtio_core_sed_record11_payload_fine_ts0)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference5 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record10_payload_address1 != main_genericstandalone_rtio_core_sed_record11_payload_address1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference5 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_134 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_135;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference6 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record12_payload_channel1 != main_genericstandalone_rtio_core_sed_record13_payload_channel1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference6 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record12_payload_fine_ts0 != main_genericstandalone_rtio_core_sed_record13_payload_fine_ts0)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference6 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record12_payload_address1 != main_genericstandalone_rtio_core_sed_record13_payload_address1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference6 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_135 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_136;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference7 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record14_payload_channel1 != main_genericstandalone_rtio_core_sed_record15_payload_channel1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference7 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record14_payload_fine_ts0 != main_genericstandalone_rtio_core_sed_record15_payload_fine_ts0)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference7 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record14_payload_address1 != main_genericstandalone_rtio_core_sed_record15_payload_address1)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference7 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_136 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_137;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference8 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record0_rec_payload_channel != main_genericstandalone_rtio_core_sed_record2_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference8 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference8 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record0_rec_payload_address != main_genericstandalone_rtio_core_sed_record2_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference8 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_137 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_138;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference9 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record1_rec_payload_channel != main_genericstandalone_rtio_core_sed_record3_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference9 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference9 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record1_rec_payload_address != main_genericstandalone_rtio_core_sed_record3_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference9 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_138 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_139;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference10 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record4_rec_payload_channel != main_genericstandalone_rtio_core_sed_record6_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference10 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference10 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record4_rec_payload_address != main_genericstandalone_rtio_core_sed_record6_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference10 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_139 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_140;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference11 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record5_rec_payload_channel != main_genericstandalone_rtio_core_sed_record7_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference11 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference11 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record5_rec_payload_address != main_genericstandalone_rtio_core_sed_record7_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference11 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_140 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_141;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference12 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record8_rec_payload_channel != main_genericstandalone_rtio_core_sed_record10_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference12 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference12 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record8_rec_payload_address != main_genericstandalone_rtio_core_sed_record10_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference12 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_141 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_142;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference13 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record9_rec_payload_channel != main_genericstandalone_rtio_core_sed_record11_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference13 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference13 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record9_rec_payload_address != main_genericstandalone_rtio_core_sed_record11_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference13 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_142 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_143;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference14 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record12_rec_payload_channel != main_genericstandalone_rtio_core_sed_record14_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference14 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference14 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record12_rec_payload_address != main_genericstandalone_rtio_core_sed_record14_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference14 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_143 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_144;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference15 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record13_rec_payload_channel != main_genericstandalone_rtio_core_sed_record15_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference15 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference15 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record13_rec_payload_address != main_genericstandalone_rtio_core_sed_record15_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference15 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_144 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_145;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference16 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record17_rec_payload_channel != main_genericstandalone_rtio_core_sed_record18_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference16 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference16 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record17_rec_payload_address != main_genericstandalone_rtio_core_sed_record18_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference16 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_145 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_146;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference17 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record21_rec_payload_channel != main_genericstandalone_rtio_core_sed_record22_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference17 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference17 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record21_rec_payload_address != main_genericstandalone_rtio_core_sed_record22_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference17 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_146 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_147;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference18 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record25_rec_payload_channel != main_genericstandalone_rtio_core_sed_record26_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference18 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference18 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record25_rec_payload_address != main_genericstandalone_rtio_core_sed_record26_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference18 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_147 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_148;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference19 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record29_rec_payload_channel != main_genericstandalone_rtio_core_sed_record30_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference19 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference19 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record29_rec_payload_address != main_genericstandalone_rtio_core_sed_record30_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference19 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_148 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_149;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference20 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record32_rec_payload_channel != main_genericstandalone_rtio_core_sed_record36_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference20 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record32_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record36_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference20 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record32_rec_payload_address != main_genericstandalone_rtio_core_sed_record36_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference20 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_149 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_150;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference21 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record33_rec_payload_channel != main_genericstandalone_rtio_core_sed_record37_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference21 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference21 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record33_rec_payload_address != main_genericstandalone_rtio_core_sed_record37_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference21 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_150 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_151;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference22 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record34_rec_payload_channel != main_genericstandalone_rtio_core_sed_record38_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference22 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference22 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record34_rec_payload_address != main_genericstandalone_rtio_core_sed_record38_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference22 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_151 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_152;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference23 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record35_rec_payload_channel != main_genericstandalone_rtio_core_sed_record39_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference23 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record35_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record39_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference23 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record35_rec_payload_address != main_genericstandalone_rtio_core_sed_record39_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference23 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_152 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_153;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference24 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record40_rec_payload_channel != main_genericstandalone_rtio_core_sed_record44_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference24 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record40_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record44_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference24 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record40_rec_payload_address != main_genericstandalone_rtio_core_sed_record44_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference24 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_153 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_154;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference25 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record41_rec_payload_channel != main_genericstandalone_rtio_core_sed_record45_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference25 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference25 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record41_rec_payload_address != main_genericstandalone_rtio_core_sed_record45_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference25 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_154 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_155;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference26 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record42_rec_payload_channel != main_genericstandalone_rtio_core_sed_record46_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference26 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference26 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record42_rec_payload_address != main_genericstandalone_rtio_core_sed_record46_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference26 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_155 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_156;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference27 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record43_rec_payload_channel != main_genericstandalone_rtio_core_sed_record47_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference27 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record43_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record47_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference27 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record43_rec_payload_address != main_genericstandalone_rtio_core_sed_record47_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference27 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_156 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_157;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference28 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record50_rec_payload_channel != main_genericstandalone_rtio_core_sed_record52_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference28 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference28 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record50_rec_payload_address != main_genericstandalone_rtio_core_sed_record52_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference28 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_157 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_158;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference29 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record51_rec_payload_channel != main_genericstandalone_rtio_core_sed_record53_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference29 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference29 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record51_rec_payload_address != main_genericstandalone_rtio_core_sed_record53_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference29 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_158 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_159;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference30 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record58_rec_payload_channel != main_genericstandalone_rtio_core_sed_record60_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference30 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference30 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record58_rec_payload_address != main_genericstandalone_rtio_core_sed_record60_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference30 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_159 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_160;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference31 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record59_rec_payload_channel != main_genericstandalone_rtio_core_sed_record61_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference31 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference31 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record59_rec_payload_address != main_genericstandalone_rtio_core_sed_record61_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference31 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_160 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_161;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference32 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record65_rec_payload_channel != main_genericstandalone_rtio_core_sed_record66_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference32 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record65_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference32 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record65_rec_payload_address != main_genericstandalone_rtio_core_sed_record66_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference32 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_161 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_162;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference33 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record67_rec_payload_channel != main_genericstandalone_rtio_core_sed_record68_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference33 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference33 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record67_rec_payload_address != main_genericstandalone_rtio_core_sed_record68_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference33 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_162 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_163;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference34 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record69_rec_payload_channel != main_genericstandalone_rtio_core_sed_record70_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference34 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record70_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference34 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record69_rec_payload_address != main_genericstandalone_rtio_core_sed_record70_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference34 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_163 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_164;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference35 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record73_rec_payload_channel != main_genericstandalone_rtio_core_sed_record74_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference35 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record73_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference35 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record73_rec_payload_address != main_genericstandalone_rtio_core_sed_record74_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference35 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_164 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_165;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference36 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record75_rec_payload_channel != main_genericstandalone_rtio_core_sed_record76_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference36 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference36 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record75_rec_payload_address != main_genericstandalone_rtio_core_sed_record76_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference36 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_165 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_166;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference37 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record77_rec_payload_channel != main_genericstandalone_rtio_core_sed_record78_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference37 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record78_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference37 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record77_rec_payload_address != main_genericstandalone_rtio_core_sed_record78_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference37 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_166 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_167;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference38 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record80_rec_payload_channel != main_genericstandalone_rtio_core_sed_record88_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference38 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record80_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record88_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference38 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record80_rec_payload_address != main_genericstandalone_rtio_core_sed_record88_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference38 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_167 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_168;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference39 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record81_rec_payload_channel != main_genericstandalone_rtio_core_sed_record89_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference39 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference39 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record81_rec_payload_address != main_genericstandalone_rtio_core_sed_record89_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference39 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_168 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_169;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference40 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record82_rec_payload_channel != main_genericstandalone_rtio_core_sed_record90_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference40 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference40 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record82_rec_payload_address != main_genericstandalone_rtio_core_sed_record90_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference40 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_169 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_170;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference41 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record83_rec_payload_channel != main_genericstandalone_rtio_core_sed_record91_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference41 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference41 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record83_rec_payload_address != main_genericstandalone_rtio_core_sed_record91_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference41 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_170 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_171;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference42 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record84_rec_payload_channel != main_genericstandalone_rtio_core_sed_record92_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference42 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference42 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record84_rec_payload_address != main_genericstandalone_rtio_core_sed_record92_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference42 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_171 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_172;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference43 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record85_rec_payload_channel != main_genericstandalone_rtio_core_sed_record93_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference43 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference43 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record85_rec_payload_address != main_genericstandalone_rtio_core_sed_record93_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference43 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_172 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_173;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference44 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record86_rec_payload_channel != main_genericstandalone_rtio_core_sed_record94_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference44 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference44 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record86_rec_payload_address != main_genericstandalone_rtio_core_sed_record94_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference44 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_173 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_174;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference45 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record87_rec_payload_channel != main_genericstandalone_rtio_core_sed_record95_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference45 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record87_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record95_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference45 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record87_rec_payload_address != main_genericstandalone_rtio_core_sed_record95_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference45 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_174 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_175;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference46 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record100_rec_payload_channel != main_genericstandalone_rtio_core_sed_record104_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference46 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference46 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record100_rec_payload_address != main_genericstandalone_rtio_core_sed_record104_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference46 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_175 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_176;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference47 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record101_rec_payload_channel != main_genericstandalone_rtio_core_sed_record105_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference47 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference47 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record101_rec_payload_address != main_genericstandalone_rtio_core_sed_record105_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference47 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_176 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_177;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference48 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record102_rec_payload_channel != main_genericstandalone_rtio_core_sed_record106_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference48 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference48 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record102_rec_payload_address != main_genericstandalone_rtio_core_sed_record106_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference48 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_177 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_178;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference49 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record103_rec_payload_channel != main_genericstandalone_rtio_core_sed_record107_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference49 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference49 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record103_rec_payload_address != main_genericstandalone_rtio_core_sed_record107_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference49 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_178 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_179;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference50 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record114_rec_payload_channel != main_genericstandalone_rtio_core_sed_record116_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference50 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record114_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference50 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record114_rec_payload_address != main_genericstandalone_rtio_core_sed_record116_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference50 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_179 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_180;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference51 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record115_rec_payload_channel != main_genericstandalone_rtio_core_sed_record117_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference51 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record115_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference51 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record115_rec_payload_address != main_genericstandalone_rtio_core_sed_record117_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference51 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_180 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_181;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference52 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record118_rec_payload_channel != main_genericstandalone_rtio_core_sed_record120_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference52 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference52 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record118_rec_payload_address != main_genericstandalone_rtio_core_sed_record120_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference52 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_181 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_182;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference53 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record119_rec_payload_channel != main_genericstandalone_rtio_core_sed_record121_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference53 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference53 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record119_rec_payload_address != main_genericstandalone_rtio_core_sed_record121_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference53 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_182 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_183;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference54 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record122_rec_payload_channel != main_genericstandalone_rtio_core_sed_record124_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference54 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record124_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference54 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record122_rec_payload_address != main_genericstandalone_rtio_core_sed_record124_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference54 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_183 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_184;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference55 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record123_rec_payload_channel != main_genericstandalone_rtio_core_sed_record125_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference55 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record125_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference55 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record123_rec_payload_address != main_genericstandalone_rtio_core_sed_record125_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference55 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_184 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_185;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference56 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record129_rec_payload_channel != main_genericstandalone_rtio_core_sed_record130_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference56 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record129_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference56 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record129_rec_payload_address != main_genericstandalone_rtio_core_sed_record130_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference56 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_185 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_186;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference57 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record131_rec_payload_channel != main_genericstandalone_rtio_core_sed_record132_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference57 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference57 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record131_rec_payload_address != main_genericstandalone_rtio_core_sed_record132_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference57 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_186 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_187;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference58 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record133_rec_payload_channel != main_genericstandalone_rtio_core_sed_record134_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference58 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference58 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record133_rec_payload_address != main_genericstandalone_rtio_core_sed_record134_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference58 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_187 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_188;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference59 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record135_rec_payload_channel != main_genericstandalone_rtio_core_sed_record136_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference59 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference59 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record135_rec_payload_address != main_genericstandalone_rtio_core_sed_record136_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference59 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_188 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_189;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference60 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record137_rec_payload_channel != main_genericstandalone_rtio_core_sed_record138_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference60 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference60 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record137_rec_payload_address != main_genericstandalone_rtio_core_sed_record138_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference60 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_189 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_190;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference61 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record139_rec_payload_channel != main_genericstandalone_rtio_core_sed_record140_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference61 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference61 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record139_rec_payload_address != main_genericstandalone_rtio_core_sed_record140_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference61 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_190 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_191;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_sed_nondata_difference62 <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record141_rec_payload_channel != main_genericstandalone_rtio_core_sed_record142_rec_payload_channel)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference62 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts != main_genericstandalone_rtio_core_sed_record142_rec_payload_fine_ts)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference62 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_sed_record141_rec_payload_address != main_genericstandalone_rtio_core_sed_record142_rec_payload_address)) begin
		main_genericstandalone_rtio_core_sed_nondata_difference62 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_191 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_din = {main_genericstandalone_rtio_core_inputcollector_record0_fifo_in_timestamp, main_genericstandalone_rtio_core_inputcollector_record0_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record0_fifo_out_timestamp, main_genericstandalone_rtio_core_inputcollector_record0_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_dout;
assign main_genericstandalone_rtio_core_inputcollector_record0_fifo_in_data = main_inout_8x0_inout_8x0_iinterface0_data;
assign main_genericstandalone_rtio_core_inputcollector_record0_fifo_in_timestamp = {main_genericstandalone_coarse_ts, main_inout_8x0_inout_8x0_iinterface0_fine_ts};
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_we = main_inout_8x0_inout_8x0_iinterface0_stb;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger0 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected0 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_re = ((main_genericstandalone_rtio_core_inputcollector_selected0 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow0));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_din = {main_genericstandalone_rtio_core_inputcollector_record1_fifo_in_timestamp, main_genericstandalone_rtio_core_inputcollector_record1_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record1_fifo_out_timestamp, main_genericstandalone_rtio_core_inputcollector_record1_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_dout;
assign main_genericstandalone_rtio_core_inputcollector_record1_fifo_in_data = main_inout_8x1_inout_8x1_iinterface1_data;
assign main_genericstandalone_rtio_core_inputcollector_record1_fifo_in_timestamp = {main_genericstandalone_coarse_ts, main_inout_8x1_inout_8x1_iinterface1_fine_ts};
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_we = main_inout_8x1_inout_8x1_iinterface1_stb;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected1 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 1'd1);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_re = ((main_genericstandalone_rtio_core_inputcollector_selected1 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow1));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_din = {main_genericstandalone_rtio_core_inputcollector_record2_fifo_in_timestamp, main_genericstandalone_rtio_core_inputcollector_record2_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record2_fifo_out_timestamp, main_genericstandalone_rtio_core_inputcollector_record2_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_dout;
assign main_genericstandalone_rtio_core_inputcollector_record2_fifo_in_data = main_inout_8x2_inout_8x2_iinterface2_data;
assign main_genericstandalone_rtio_core_inputcollector_record2_fifo_in_timestamp = {main_genericstandalone_coarse_ts, main_inout_8x2_inout_8x2_iinterface2_fine_ts};
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_we = main_inout_8x2_inout_8x2_iinterface2_stb;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger2 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected2 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 2'd2);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_re = ((main_genericstandalone_rtio_core_inputcollector_selected2 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow2));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_din = {main_genericstandalone_rtio_core_inputcollector_record3_fifo_in_timestamp, main_genericstandalone_rtio_core_inputcollector_record3_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record3_fifo_out_timestamp, main_genericstandalone_rtio_core_inputcollector_record3_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_dout;
assign main_genericstandalone_rtio_core_inputcollector_record3_fifo_in_data = main_inout_8x3_inout_8x3_iinterface3_data;
assign main_genericstandalone_rtio_core_inputcollector_record3_fifo_in_timestamp = {main_genericstandalone_coarse_ts, main_inout_8x3_inout_8x3_iinterface3_fine_ts};
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_we = main_inout_8x3_inout_8x3_iinterface3_stb;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger3 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected3 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 2'd3);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_re = ((main_genericstandalone_rtio_core_inputcollector_selected3 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow3));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_din = {main_genericstandalone_rtio_core_inputcollector_record4_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record4_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_dout;
assign main_genericstandalone_rtio_core_inputcollector_record4_fifo_in_data = main_spimaster0_iinterface0_data0;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_we = main_spimaster0_iinterface0_stb0;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger4 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected4 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 5'd16);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_re = ((main_genericstandalone_rtio_core_inputcollector_selected4 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow4));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_din = {main_genericstandalone_rtio_core_inputcollector_record5_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record5_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_dout;
assign main_genericstandalone_rtio_core_inputcollector_record5_fifo_in_data = main_spimaster1_iinterface1_data0;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_we = main_spimaster1_iinterface1_stb0;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger5 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected5 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 5'd22);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_re = ((main_genericstandalone_rtio_core_inputcollector_selected5 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow5));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_din = {main_genericstandalone_rtio_core_inputcollector_record6_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record6_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_dout;
assign main_genericstandalone_rtio_core_inputcollector_record6_fifo_in_data = main_spimaster0_iinterface0_data1;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_we = main_spimaster0_iinterface0_stb1;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger6 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected6 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 5'd28);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_re = ((main_genericstandalone_rtio_core_inputcollector_selected6 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow6));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_din = {main_genericstandalone_rtio_core_inputcollector_record7_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record7_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_dout;
assign main_genericstandalone_rtio_core_inputcollector_record7_fifo_in_data = main_spimaster1_iinterface1_data1;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_we = main_spimaster1_iinterface1_stb1;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger7 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected7 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 5'd29);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_re = ((main_genericstandalone_rtio_core_inputcollector_selected7 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow7));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_din = {main_genericstandalone_rtio_core_inputcollector_record8_fifo_in_data};
assign {main_genericstandalone_rtio_core_inputcollector_record8_fifo_out_data} = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_dout;
assign main_genericstandalone_rtio_core_inputcollector_record8_fifo_in_data = main_spimaster2_iinterface2_data;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_we = main_spimaster2_iinterface2_stb;
assign main_genericstandalone_rtio_core_inputcollector_overflow_trigger8 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_we & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_writable));
assign main_genericstandalone_rtio_core_inputcollector_selected8 = (main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 5'd31);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_re = ((main_genericstandalone_rtio_core_inputcollector_selected8 & main_genericstandalone_rtio_core_inputcollector_i_ack) & (~main_genericstandalone_rtio_core_inputcollector_overflow8));
assign main_genericstandalone_rtio_core_inputcollector_i_status_raw = builder_comb_rhs_self10;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_readable);

// synthesis translate_off
reg dummy_d_192;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_adr <= 6'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_produce;
	end
// synthesis translate_off
	dummy_d_192 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 != 7'd64);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 != 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_readable);

// synthesis translate_off
reg dummy_d_193;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_adr <= 6'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_produce;
	end
// synthesis translate_off
	dummy_d_193 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 != 7'd64);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 != 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_readable);

// synthesis translate_off
reg dummy_d_194;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_adr <= 6'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_produce;
	end
// synthesis translate_off
	dummy_d_194 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 != 7'd64);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 != 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_readable);

// synthesis translate_off
reg dummy_d_195;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_adr <= 6'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_produce;
	end
// synthesis translate_off
	dummy_d_195 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 != 7'd64);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 != 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_readable);

// synthesis translate_off
reg dummy_d_196;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_adr <= 2'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_produce;
	end
// synthesis translate_off
	dummy_d_196 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 != 3'd4);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 != 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_readable);

// synthesis translate_off
reg dummy_d_197;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_adr <= 2'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_produce;
	end
// synthesis translate_off
	dummy_d_197 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 != 3'd4);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 != 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_readable);

// synthesis translate_off
reg dummy_d_198;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_adr <= 2'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_produce;
	end
// synthesis translate_off
	dummy_d_198 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 != 3'd4);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 != 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_readable);

// synthesis translate_off
reg dummy_d_199;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_adr <= 2'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_produce;
	end
// synthesis translate_off
	dummy_d_199 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 != 3'd4);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 != 1'd0);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_re = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_readable & ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_readable) | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_re));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level1 = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 + main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_readable);

// synthesis translate_off
reg dummy_d_200;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_adr <= 2'd0;
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_replace) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_adr <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_adr <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_produce;
	end
// synthesis translate_off
	dummy_d_200 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_dat_w = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_din;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_we = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_we & (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_writable | main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_replace));
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_do_read = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_readable & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_re);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_adr = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_consume;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_dout = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_dat_r;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_re = main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_do_read;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_writable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 != 3'd4);
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_readable = (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 != 1'd0);
assign main_genericstandalone_rtio_core_o_collision_sync_ps_i = (main_genericstandalone_rtio_core_o_collision_sync_i & (~main_genericstandalone_rtio_core_o_collision_sync_blind));
assign main_genericstandalone_rtio_core_o_collision_sync_ps_ack_i = main_genericstandalone_rtio_core_o_collision_sync_ps_o;
assign main_genericstandalone_rtio_core_o_collision_sync_o = main_genericstandalone_rtio_core_o_collision_sync_ps_o;
assign main_genericstandalone_rtio_core_o_collision_sync_ps_o = (main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_o ^ main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_o_r);
assign main_genericstandalone_rtio_core_o_collision_sync_ps_ack_o = (main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_o ^ main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_o_r);
assign main_genericstandalone_rtio_core_o_busy_sync_ps_i = (main_genericstandalone_rtio_core_o_busy_sync_i & (~main_genericstandalone_rtio_core_o_busy_sync_blind));
assign main_genericstandalone_rtio_core_o_busy_sync_ps_ack_i = main_genericstandalone_rtio_core_o_busy_sync_ps_o;
assign main_genericstandalone_rtio_core_o_busy_sync_o = main_genericstandalone_rtio_core_o_busy_sync_ps_o;
assign main_genericstandalone_rtio_core_o_busy_sync_ps_o = (main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_o ^ main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_o_r);
assign main_genericstandalone_rtio_core_o_busy_sync_ps_ack_o = (main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_o ^ main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_o_r);
assign main_genericstandalone_rtio_now_hi_w = main_genericstandalone_rtio_now[63:32];
assign main_genericstandalone_rtio_now_lo_w = main_genericstandalone_rtio_now[31:0];

// synthesis translate_off
reg dummy_d_201;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_cri_cmd <= 2'd0;
	main_genericstandalone_rtio_cri_cmd <= 1'd0;
	if (main_genericstandalone_rtio_o_data_re) begin
		main_genericstandalone_rtio_cri_cmd <= 1'd1;
	end
	if (main_genericstandalone_rtio_i_timeout_re) begin
		main_genericstandalone_rtio_cri_cmd <= 2'd2;
	end
// synthesis translate_off
	dummy_d_201 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_cri_chan_sel = main_genericstandalone_rtio_target_storage[31:8];
assign main_genericstandalone_rtio_cri_o_timestamp = main_genericstandalone_rtio_now;
assign main_genericstandalone_rtio_cri_o_data = main_genericstandalone_rtio_o_data_storage;
assign main_genericstandalone_rtio_cri_o_address = main_genericstandalone_rtio_target_storage[7:0];
assign main_genericstandalone_rtio_o_status_status = main_genericstandalone_rtio_cri_o_status;
assign main_genericstandalone_rtio_cri_i_timeout = main_genericstandalone_rtio_i_timeout_storage;
assign main_genericstandalone_rtio_i_data_status = main_genericstandalone_rtio_cri_i_data;
assign main_genericstandalone_rtio_i_timestamp_status = main_genericstandalone_rtio_cri_i_timestamp;
assign main_genericstandalone_rtio_i_status_status = main_genericstandalone_rtio_cri_i_status;
assign main_genericstandalone_rtio_o_data_dat_w = 1'd0;
assign main_genericstandalone_rtio_o_data_we = main_genericstandalone_rtio_target_re;
assign main_genericstandalone_dma_fifo_sink_stb = main_genericstandalone_dma_dma_source_stb;
assign main_genericstandalone_dma_dma_source_ack = main_genericstandalone_dma_fifo_sink_ack;
assign main_genericstandalone_dma_fifo_sink_last = main_genericstandalone_dma_dma_source_last;
assign main_genericstandalone_dma_fifo_sink_eop = main_genericstandalone_dma_dma_source_eop;
assign main_genericstandalone_dma_fifo_sink_payload_data = main_genericstandalone_dma_dma_source_payload_data;
assign main_genericstandalone_dma_rawslicer_sink_stb = main_genericstandalone_dma_fifo_source_stb;
assign main_genericstandalone_dma_fifo_source_ack = main_genericstandalone_dma_rawslicer_sink_ack;
assign main_genericstandalone_dma_rawslicer_sink_last = main_genericstandalone_dma_fifo_source_last;
assign main_genericstandalone_dma_rawslicer_sink_eop = main_genericstandalone_dma_fifo_source_eop;
assign main_genericstandalone_dma_rawslicer_sink_payload_data = main_genericstandalone_dma_fifo_source_payload_data;
assign main_genericstandalone_dma_time_offset_sink_stb = main_genericstandalone_dma_record_converter_source_stb;
assign main_genericstandalone_dma_record_converter_source_ack = main_genericstandalone_dma_time_offset_sink_ack;
assign main_genericstandalone_dma_time_offset_sink_last = main_genericstandalone_dma_record_converter_source_last;
assign main_genericstandalone_dma_time_offset_sink_eop = main_genericstandalone_dma_record_converter_source_eop;
assign main_genericstandalone_dma_time_offset_sink_payload_length = main_genericstandalone_dma_record_converter_source_payload_length;
assign main_genericstandalone_dma_time_offset_sink_payload_channel = main_genericstandalone_dma_record_converter_source_payload_channel;
assign main_genericstandalone_dma_time_offset_sink_payload_timestamp = main_genericstandalone_dma_record_converter_source_payload_timestamp;
assign main_genericstandalone_dma_time_offset_sink_payload_address = main_genericstandalone_dma_record_converter_source_payload_address;
assign main_genericstandalone_dma_time_offset_sink_payload_data = main_genericstandalone_dma_record_converter_source_payload_data;
assign main_genericstandalone_dma_cri_master_sink_stb = main_genericstandalone_dma_time_offset_source_stb;
assign main_genericstandalone_dma_time_offset_source_ack = main_genericstandalone_dma_cri_master_sink_ack;
assign main_genericstandalone_dma_cri_master_sink_last = main_genericstandalone_dma_time_offset_source_last;
assign main_genericstandalone_dma_cri_master_sink_eop = main_genericstandalone_dma_time_offset_source_eop;
assign main_genericstandalone_dma_cri_master_sink_payload_length = main_genericstandalone_dma_time_offset_source_payload_length;
assign main_genericstandalone_dma_cri_master_sink_payload_channel = main_genericstandalone_dma_time_offset_source_payload_channel;
assign main_genericstandalone_dma_cri_master_sink_payload_timestamp = main_genericstandalone_dma_time_offset_source_payload_timestamp;
assign main_genericstandalone_dma_cri_master_sink_payload_address = main_genericstandalone_dma_time_offset_source_payload_address;
assign main_genericstandalone_dma_cri_master_sink_payload_data = main_genericstandalone_dma_time_offset_source_payload_data;
assign main_genericstandalone_dma_dma_bus_stb = (main_genericstandalone_dma_dma_sink_stb & main_genericstandalone_dma_dma_source_ack);
assign main_genericstandalone_dma_dma_last = (main_genericstandalone_dma_dma_transfer_cyc == 1'd0);
assign main_genericstandalone_dma_dma_transfer_cyc_rst = ((main_genericstandalone_dma_dma_source_stb & main_genericstandalone_dma_dma_source_ack) & (main_genericstandalone_dma_dma_sink_eop | main_genericstandalone_dma_dma_last));
assign main_genericstandalone_dma_dma_transfer_cyc_ce = (main_genericstandalone_dma_dma_source_stb & main_genericstandalone_dma_dma_source_ack);
assign main_genericstandalone_interface0_bus_cyc = main_genericstandalone_dma_dma_bus_stb;
assign main_genericstandalone_interface0_bus_stb = main_genericstandalone_dma_dma_bus_stb;
assign main_genericstandalone_interface0_bus_cti = ((main_genericstandalone_dma_dma_sink_eop | main_genericstandalone_dma_dma_last) ? 3'd7 : 2'd2);
assign main_genericstandalone_interface0_bus_adr = main_genericstandalone_dma_dma_sink_payload_address;
assign main_genericstandalone_dma_dma_sink_ack = main_genericstandalone_interface0_bus_ack;
assign main_genericstandalone_dma_dma_source_stb = main_genericstandalone_interface0_bus_ack;
assign main_genericstandalone_dma_dma_source_payload_data = {{builder_slice_proxy15[7:0], builder_slice_proxy14[15:8], builder_slice_proxy13[23:16], builder_slice_proxy12[31:24], builder_slice_proxy11[39:32], builder_slice_proxy10[47:40], builder_slice_proxy9[55:48], builder_slice_proxy8[63:56]}, {builder_slice_proxy7[7:0], builder_slice_proxy6[15:8], builder_slice_proxy5[23:16], builder_slice_proxy4[31:24], builder_slice_proxy3[39:32], builder_slice_proxy2[47:40], builder_slice_proxy1[55:48], builder_slice_proxy0[63:56]}};
assign main_genericstandalone_dma_dma_source_last = (main_genericstandalone_dma_dma_sink_eop | main_genericstandalone_dma_dma_last);
assign main_genericstandalone_dma_dma_source_eop = main_genericstandalone_dma_dma_sink_eop;
assign main_genericstandalone_dma_fifo_syncfifo_din = {main_genericstandalone_dma_fifo_fifo_in_eop, main_genericstandalone_dma_fifo_fifo_in_payload_data};
assign {main_genericstandalone_dma_fifo_fifo_out_eop, main_genericstandalone_dma_fifo_fifo_out_payload_data} = main_genericstandalone_dma_fifo_syncfifo_dout;
assign main_genericstandalone_dma_fifo_fifo_in_eop = main_genericstandalone_dma_fifo_sink_eop;
assign main_genericstandalone_dma_fifo_fifo_in_payload_data = main_genericstandalone_dma_fifo_sink_payload_data;
assign main_genericstandalone_dma_fifo_source_stb = main_genericstandalone_dma_fifo_readable;
assign main_genericstandalone_dma_fifo_source_eop = main_genericstandalone_dma_fifo_fifo_out_eop;
assign main_genericstandalone_dma_fifo_source_payload_data = main_genericstandalone_dma_fifo_fifo_out_payload_data;
assign main_genericstandalone_dma_fifo_re = main_genericstandalone_dma_fifo_source_ack;
assign main_genericstandalone_dma_fifo_do_write = (main_genericstandalone_dma_fifo_syncfifo_we & main_genericstandalone_dma_fifo_syncfifo_writable);

// synthesis translate_off
reg dummy_d_202;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_dma_fifo_syncfifo_we <= 1'd0;
	main_genericstandalone_dma_fifo_syncfifo_we <= main_genericstandalone_dma_fifo_sink_stb;
	main_genericstandalone_dma_fifo_syncfifo_we <= (main_genericstandalone_dma_fifo_sink_stb & main_genericstandalone_dma_fifo_sink_ack);
// synthesis translate_off
	dummy_d_202 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_203;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_dma_fifo_sink_ack <= 1'd0;
	main_genericstandalone_dma_fifo_sink_ack <= main_genericstandalone_dma_fifo_syncfifo_writable;
	main_genericstandalone_dma_fifo_sink_ack <= (main_genericstandalone_dma_fifo_syncfifo_writable & (main_genericstandalone_dma_fifo_almost_empty | main_genericstandalone_dma_fifo_recv_activated));
// synthesis translate_off
	dummy_d_203 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_dma_fifo_syncfifo_re = (main_genericstandalone_dma_fifo_syncfifo_readable & ((~main_genericstandalone_dma_fifo_readable) | main_genericstandalone_dma_fifo_re));
assign main_genericstandalone_dma_fifo_level1 = (main_genericstandalone_dma_fifo_level0 + main_genericstandalone_dma_fifo_readable);
assign main_genericstandalone_dma_fifo_almost_empty = (main_genericstandalone_dma_fifo_level1 <= 7'd64);

// synthesis translate_off
reg dummy_d_204;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_dma_fifo_wrport_adr <= 7'd0;
	if (main_genericstandalone_dma_fifo_replace) begin
		main_genericstandalone_dma_fifo_wrport_adr <= (main_genericstandalone_dma_fifo_produce - 1'd1);
	end else begin
		main_genericstandalone_dma_fifo_wrport_adr <= main_genericstandalone_dma_fifo_produce;
	end
// synthesis translate_off
	dummy_d_204 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_dma_fifo_wrport_dat_w = main_genericstandalone_dma_fifo_syncfifo_din;
assign main_genericstandalone_dma_fifo_wrport_we = (main_genericstandalone_dma_fifo_syncfifo_we & (main_genericstandalone_dma_fifo_syncfifo_writable | main_genericstandalone_dma_fifo_replace));
assign main_genericstandalone_dma_fifo_do_read = (main_genericstandalone_dma_fifo_syncfifo_readable & main_genericstandalone_dma_fifo_syncfifo_re);
assign main_genericstandalone_dma_fifo_rdport_adr = main_genericstandalone_dma_fifo_consume;
assign main_genericstandalone_dma_fifo_syncfifo_dout = main_genericstandalone_dma_fifo_rdport_dat_r;
assign main_genericstandalone_dma_fifo_rdport_re = main_genericstandalone_dma_fifo_do_read;
assign main_genericstandalone_dma_fifo_syncfifo_writable = (main_genericstandalone_dma_fifo_level0 != 8'd128);
assign main_genericstandalone_dma_fifo_syncfifo_readable = (main_genericstandalone_dma_fifo_level0 != 1'd0);
assign main_genericstandalone_dma_rawslicer_source = main_genericstandalone_dma_rawslicer_buf[615:0];

// synthesis translate_off
reg dummy_d_205;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_dma_rawslicer_sink_ack <= 1'd0;
	main_genericstandalone_dma_rawslicer_source_stb <= 1'd0;
	main_genericstandalone_dma_rawslicer_flush_done <= 1'd0;
	main_genericstandalone_dma_rawslicer_next_level <= 7'd0;
	main_genericstandalone_dma_rawslicer_load_buf <= 1'd0;
	main_genericstandalone_dma_rawslicer_shift_buf <= 1'd0;
	builder_clockdomainsrenamer_resetinserter_next_state <= 2'd0;
	main_genericstandalone_dma_rawslicer_next_level <= main_genericstandalone_dma_rawslicer_level;
	builder_clockdomainsrenamer_resetinserter_next_state <= builder_clockdomainsrenamer_resetinserter_state;
	case (builder_clockdomainsrenamer_resetinserter_state)
		1'd1: begin
			main_genericstandalone_dma_rawslicer_source_stb <= 1'd1;
			main_genericstandalone_dma_rawslicer_shift_buf <= 1'd1;
			main_genericstandalone_dma_rawslicer_next_level <= (main_genericstandalone_dma_rawslicer_level - main_genericstandalone_dma_rawslicer_source_consume);
			if ((main_genericstandalone_dma_rawslicer_next_level < 7'd77)) begin
				builder_clockdomainsrenamer_resetinserter_next_state <= 1'd0;
			end
			if (main_genericstandalone_dma_rawslicer_flush) begin
				builder_clockdomainsrenamer_resetinserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_genericstandalone_dma_rawslicer_next_level <= 1'd0;
			main_genericstandalone_dma_rawslicer_sink_ack <= 1'd1;
			if ((main_genericstandalone_dma_rawslicer_sink_stb & main_genericstandalone_dma_rawslicer_sink_eop)) begin
				main_genericstandalone_dma_rawslicer_flush_done <= 1'd1;
				builder_clockdomainsrenamer_resetinserter_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_dma_rawslicer_sink_ack <= 1'd1;
			main_genericstandalone_dma_rawslicer_load_buf <= 1'd1;
			if (main_genericstandalone_dma_rawslicer_sink_stb) begin
				main_genericstandalone_dma_rawslicer_next_level <= (main_genericstandalone_dma_rawslicer_level + 5'd16);
			end
			if ((main_genericstandalone_dma_rawslicer_next_level >= 7'd77)) begin
				builder_clockdomainsrenamer_resetinserter_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_205 <= dummy_s;
// synthesis translate_on
end
assign {main_genericstandalone_dma_record_converter_record_raw_data, main_genericstandalone_dma_record_converter_record_raw_address, main_genericstandalone_dma_record_converter_record_raw_timestamp, main_genericstandalone_dma_record_converter_record_raw_channel, main_genericstandalone_dma_record_converter_record_raw_length} = main_genericstandalone_dma_rawslicer_source;
assign main_genericstandalone_dma_record_converter_source_payload_channel = main_genericstandalone_dma_record_converter_record_raw_channel;
assign main_genericstandalone_dma_record_converter_source_payload_timestamp = main_genericstandalone_dma_record_converter_record_raw_timestamp;
assign main_genericstandalone_dma_record_converter_source_payload_address = main_genericstandalone_dma_record_converter_record_raw_address;

// synthesis translate_off
reg dummy_d_206;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_dma_record_converter_source_payload_data <= 512'd0;
	case (main_genericstandalone_dma_record_converter_record_raw_length)
		4'd14: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[7:0];
		end
		4'd15: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[15:0];
		end
		5'd16: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[23:0];
		end
		5'd17: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[31:0];
		end
		5'd18: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[39:0];
		end
		5'd19: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[47:0];
		end
		5'd20: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[55:0];
		end
		5'd21: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[63:0];
		end
		5'd22: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[71:0];
		end
		5'd23: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[79:0];
		end
		5'd24: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[87:0];
		end
		5'd25: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[95:0];
		end
		5'd26: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[103:0];
		end
		5'd27: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[111:0];
		end
		5'd28: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[119:0];
		end
		5'd29: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[127:0];
		end
		5'd30: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[135:0];
		end
		5'd31: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[143:0];
		end
		6'd32: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[151:0];
		end
		6'd33: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[159:0];
		end
		6'd34: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[167:0];
		end
		6'd35: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[175:0];
		end
		6'd36: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[183:0];
		end
		6'd37: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[191:0];
		end
		6'd38: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[199:0];
		end
		6'd39: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[207:0];
		end
		6'd40: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[215:0];
		end
		6'd41: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[223:0];
		end
		6'd42: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[231:0];
		end
		6'd43: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[239:0];
		end
		6'd44: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[247:0];
		end
		6'd45: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[255:0];
		end
		6'd46: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[263:0];
		end
		6'd47: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[271:0];
		end
		6'd48: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[279:0];
		end
		6'd49: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[287:0];
		end
		6'd50: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[295:0];
		end
		6'd51: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[303:0];
		end
		6'd52: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[311:0];
		end
		6'd53: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[319:0];
		end
		6'd54: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[327:0];
		end
		6'd55: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[335:0];
		end
		6'd56: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[343:0];
		end
		6'd57: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[351:0];
		end
		6'd58: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[359:0];
		end
		6'd59: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[367:0];
		end
		6'd60: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[375:0];
		end
		6'd61: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[383:0];
		end
		6'd62: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[391:0];
		end
		6'd63: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[399:0];
		end
		7'd64: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[407:0];
		end
		7'd65: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[415:0];
		end
		7'd66: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[423:0];
		end
		7'd67: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[431:0];
		end
		7'd68: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[439:0];
		end
		7'd69: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[447:0];
		end
		7'd70: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[455:0];
		end
		7'd71: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[463:0];
		end
		7'd72: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[471:0];
		end
		7'd73: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[479:0];
		end
		7'd74: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[487:0];
		end
		7'd75: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[495:0];
		end
		7'd76: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[503:0];
		end
		7'd77: begin
			main_genericstandalone_dma_record_converter_source_payload_data <= main_genericstandalone_dma_record_converter_record_raw_data[511:0];
		end
	endcase
// synthesis translate_off
	dummy_d_206 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_207;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_dma_rawslicer_source_consume <= 7'd0;
	main_genericstandalone_dma_rawslicer_flush <= 1'd0;
	main_genericstandalone_dma_record_converter_source_stb <= 1'd0;
	main_genericstandalone_dma_record_converter_source_eop <= 1'd0;
	main_genericstandalone_dma_record_converter_end_marker_found <= 1'd0;
	builder_clockdomainsrenamer_recordconverter_next_state <= 2'd0;
	builder_clockdomainsrenamer_recordconverter_next_state <= builder_clockdomainsrenamer_recordconverter_state;
	case (builder_clockdomainsrenamer_recordconverter_state)
		1'd1: begin
			main_genericstandalone_dma_record_converter_end_marker_found <= 1'd1;
			if (main_genericstandalone_dma_record_converter_flush) begin
				main_genericstandalone_dma_rawslicer_flush <= 1'd1;
				builder_clockdomainsrenamer_recordconverter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (main_genericstandalone_dma_rawslicer_flush_done) begin
				builder_clockdomainsrenamer_recordconverter_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_genericstandalone_dma_record_converter_source_eop <= 1'd1;
			main_genericstandalone_dma_record_converter_source_stb <= 1'd1;
			if (main_genericstandalone_dma_record_converter_source_ack) begin
				builder_clockdomainsrenamer_recordconverter_next_state <= 1'd0;
			end
		end
		default: begin
			if (main_genericstandalone_dma_rawslicer_source_stb) begin
				if ((main_genericstandalone_dma_record_converter_record_raw_length == 1'd0)) begin
					builder_clockdomainsrenamer_recordconverter_next_state <= 1'd1;
				end else begin
					main_genericstandalone_dma_record_converter_source_stb <= 1'd1;
				end
			end
			if (main_genericstandalone_dma_record_converter_source_ack) begin
				main_genericstandalone_dma_rawslicer_source_consume <= main_genericstandalone_dma_record_converter_record_raw_length;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_207 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_dma_time_offset_sink_ack = (~main_genericstandalone_dma_time_offset_source_stb);
assign main_genericstandalone_dma_cri_master_cri_chan_sel = main_genericstandalone_dma_cri_master_sink_payload_channel;
assign main_genericstandalone_dma_cri_master_cri_o_timestamp = main_genericstandalone_dma_cri_master_sink_payload_timestamp;
assign main_genericstandalone_dma_cri_master_cri_o_address = main_genericstandalone_dma_cri_master_sink_payload_address;
assign main_genericstandalone_dma_cri_master_cri_o_data = main_genericstandalone_dma_cri_master_sink_payload_data;

// synthesis translate_off
reg dummy_d_208;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_dma_cri_master_sink_ack <= 1'd0;
	main_genericstandalone_dma_cri_master_cri_cmd <= 2'd0;
	main_genericstandalone_dma_cri_master_busy <= 1'd0;
	main_genericstandalone_dma_cri_master_underflow_trigger <= 1'd0;
	main_genericstandalone_dma_cri_master_link_error_trigger <= 1'd0;
	builder_clockdomainsrenamer_crimaster_next_state <= 3'd0;
	builder_clockdomainsrenamer_crimaster_next_state <= builder_clockdomainsrenamer_crimaster_state;
	case (builder_clockdomainsrenamer_crimaster_state)
		1'd1: begin
			main_genericstandalone_dma_cri_master_busy <= 1'd1;
			main_genericstandalone_dma_cri_master_cri_cmd <= 1'd1;
			builder_clockdomainsrenamer_crimaster_next_state <= 2'd2;
		end
		2'd2: begin
			main_genericstandalone_dma_cri_master_busy <= 1'd1;
			if ((main_genericstandalone_dma_cri_master_cri_o_status == 1'd0)) begin
				main_genericstandalone_dma_cri_master_sink_ack <= 1'd1;
				builder_clockdomainsrenamer_crimaster_next_state <= 1'd0;
			end
			if (main_genericstandalone_dma_cri_master_cri_o_status[1]) begin
				builder_clockdomainsrenamer_crimaster_next_state <= 2'd3;
			end
			if (main_genericstandalone_dma_cri_master_cri_o_status[2]) begin
				builder_clockdomainsrenamer_crimaster_next_state <= 3'd4;
			end
		end
		2'd3: begin
			main_genericstandalone_dma_cri_master_busy <= 1'd1;
			main_genericstandalone_dma_cri_master_underflow_trigger <= 1'd1;
			main_genericstandalone_dma_cri_master_sink_ack <= 1'd1;
			builder_clockdomainsrenamer_crimaster_next_state <= 1'd0;
		end
		3'd4: begin
			main_genericstandalone_dma_cri_master_busy <= 1'd1;
			main_genericstandalone_dma_cri_master_link_error_trigger <= 1'd1;
			main_genericstandalone_dma_cri_master_sink_ack <= 1'd1;
			builder_clockdomainsrenamer_crimaster_next_state <= 1'd0;
		end
		default: begin
			if ((main_genericstandalone_dma_cri_master_error_w == 1'd0)) begin
				if (main_genericstandalone_dma_cri_master_sink_stb) begin
					if (main_genericstandalone_dma_cri_master_sink_eop) begin
						main_genericstandalone_dma_cri_master_sink_ack <= 1'd1;
					end else begin
						builder_clockdomainsrenamer_crimaster_next_state <= 1'd1;
					end
				end
			end else begin
				main_genericstandalone_dma_cri_master_sink_ack <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_208 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_209;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_dma_enable_enable_w <= 1'd0;
	main_genericstandalone_dma_flow_enable <= 1'd0;
	main_genericstandalone_dma_record_converter_flush <= 1'd0;
	builder_clockdomainsrenamer_fsm_next_state <= 3'd0;
	builder_clockdomainsrenamer_fsm_next_state <= builder_clockdomainsrenamer_fsm_state;
	case (builder_clockdomainsrenamer_fsm_state)
		1'd1: begin
			main_genericstandalone_dma_enable_enable_w <= 1'd1;
			main_genericstandalone_dma_flow_enable <= 1'd1;
			if (main_genericstandalone_dma_record_converter_end_marker_found) begin
				builder_clockdomainsrenamer_fsm_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_genericstandalone_dma_enable_enable_w <= 1'd1;
			main_genericstandalone_dma_record_converter_flush <= 1'd1;
			builder_clockdomainsrenamer_fsm_next_state <= 2'd3;
		end
		2'd3: begin
			main_genericstandalone_dma_enable_enable_w <= 1'd1;
			if (((main_genericstandalone_dma_cri_master_sink_stb & main_genericstandalone_dma_cri_master_sink_ack) & main_genericstandalone_dma_cri_master_sink_eop)) begin
				builder_clockdomainsrenamer_fsm_next_state <= 3'd4;
			end
		end
		3'd4: begin
			main_genericstandalone_dma_enable_enable_w <= 1'd1;
			if ((~main_genericstandalone_dma_cri_master_busy)) begin
				builder_clockdomainsrenamer_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			if (main_genericstandalone_dma_enable_enable_re) begin
				builder_clockdomainsrenamer_fsm_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_209 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_target0_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_target0_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 1'd0));
assign main_genericstandalone_rtio_now_hi_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_rtio_now_hi_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 1'd1));
assign main_genericstandalone_rtio_now_lo_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_rtio_now_lo_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 2'd2));
assign main_genericstandalone_o_data15_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data15_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 2'd3));
assign main_genericstandalone_o_data14_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data14_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 3'd4));
assign main_genericstandalone_o_data13_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data13_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 3'd5));
assign main_genericstandalone_o_data12_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data12_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 3'd6));
assign main_genericstandalone_o_data11_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data11_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 3'd7));
assign main_genericstandalone_o_data10_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data10_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 4'd8));
assign main_genericstandalone_o_data9_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data9_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 4'd9));
assign main_genericstandalone_o_data8_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data8_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 4'd10));
assign main_genericstandalone_o_data7_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data7_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 4'd11));
assign main_genericstandalone_o_data6_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data6_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 4'd12));
assign main_genericstandalone_o_data5_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data5_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 4'd13));
assign main_genericstandalone_o_data4_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data4_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 4'd14));
assign main_genericstandalone_o_data3_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data3_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 4'd15));
assign main_genericstandalone_o_data2_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data2_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd16));
assign main_genericstandalone_o_data1_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data1_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd17));
assign main_genericstandalone_o_data0_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_o_data0_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd18));
assign main_genericstandalone_o_status_r = main_genericstandalone_interface0_csr_bus_dat_w[2:0];
assign main_genericstandalone_o_status_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd19));
assign main_genericstandalone_i_timeout1_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_i_timeout1_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd20));
assign main_genericstandalone_i_timeout0_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_i_timeout0_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd21));
assign main_genericstandalone_i_data_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_i_data_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd22));
assign main_genericstandalone_i_timestamp1_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_i_timestamp1_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd23));
assign main_genericstandalone_i_timestamp0_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_i_timestamp0_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd24));
assign main_genericstandalone_i_status_r = main_genericstandalone_interface0_csr_bus_dat_w[3:0];
assign main_genericstandalone_i_status_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd25));
assign main_genericstandalone_counter1_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_counter1_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd26));
assign main_genericstandalone_counter0_r = main_genericstandalone_interface0_csr_bus_dat_w[31:0];
assign main_genericstandalone_counter0_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd27));
assign main_genericstandalone_rtio_counter_update_r = main_genericstandalone_interface0_csr_bus_dat_w[0];
assign main_genericstandalone_rtio_counter_update_re = ((((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb) & (~main_genericstandalone_interface0_csr_bus_ack)) & main_genericstandalone_interface0_csr_bus_we) & (main_genericstandalone_interface0_csr_bus_adr[4:0] == 5'd28));
assign main_genericstandalone_rtio_target_storage = main_genericstandalone_rtio_target_storage_full[31:0];
assign main_genericstandalone_target0_w = main_genericstandalone_rtio_target_storage_full[31:0];
assign main_genericstandalone_rtio_o_data_storage = main_genericstandalone_rtio_o_data_storage_full[511:0];
assign main_genericstandalone_o_data15_w = main_genericstandalone_rtio_o_data_storage_full[511:480];
assign main_genericstandalone_o_data14_w = main_genericstandalone_rtio_o_data_storage_full[479:448];
assign main_genericstandalone_o_data13_w = main_genericstandalone_rtio_o_data_storage_full[447:416];
assign main_genericstandalone_o_data12_w = main_genericstandalone_rtio_o_data_storage_full[415:384];
assign main_genericstandalone_o_data11_w = main_genericstandalone_rtio_o_data_storage_full[383:352];
assign main_genericstandalone_o_data10_w = main_genericstandalone_rtio_o_data_storage_full[351:320];
assign main_genericstandalone_o_data9_w = main_genericstandalone_rtio_o_data_storage_full[319:288];
assign main_genericstandalone_o_data8_w = main_genericstandalone_rtio_o_data_storage_full[287:256];
assign main_genericstandalone_o_data7_w = main_genericstandalone_rtio_o_data_storage_full[255:224];
assign main_genericstandalone_o_data6_w = main_genericstandalone_rtio_o_data_storage_full[223:192];
assign main_genericstandalone_o_data5_w = main_genericstandalone_rtio_o_data_storage_full[191:160];
assign main_genericstandalone_o_data4_w = main_genericstandalone_rtio_o_data_storage_full[159:128];
assign main_genericstandalone_o_data3_w = main_genericstandalone_rtio_o_data_storage_full[127:96];
assign main_genericstandalone_o_data2_w = main_genericstandalone_rtio_o_data_storage_full[95:64];
assign main_genericstandalone_o_data1_w = main_genericstandalone_rtio_o_data_storage_full[63:32];
assign main_genericstandalone_o_data0_w = main_genericstandalone_rtio_o_data_storage_full[31:0];
assign main_genericstandalone_o_status_w = main_genericstandalone_rtio_o_status_status[2:0];
assign main_genericstandalone_rtio_i_timeout_storage = main_genericstandalone_rtio_i_timeout_storage_full[63:0];
assign main_genericstandalone_i_timeout1_w = main_genericstandalone_rtio_i_timeout_storage_full[63:32];
assign main_genericstandalone_i_timeout0_w = main_genericstandalone_rtio_i_timeout_storage_full[31:0];
assign main_genericstandalone_i_data_w = main_genericstandalone_rtio_i_data_status[31:0];
assign main_genericstandalone_i_timestamp1_w = main_genericstandalone_rtio_i_timestamp_status[63:32];
assign main_genericstandalone_i_timestamp0_w = main_genericstandalone_rtio_i_timestamp_status[31:0];
assign main_genericstandalone_i_status_w = main_genericstandalone_rtio_i_status_status[3:0];
assign main_genericstandalone_counter1_w = main_genericstandalone_rtio_counter_status[63:32];
assign main_genericstandalone_counter0_w = main_genericstandalone_rtio_counter_status[31:0];
assign main_genericstandalone_dma_enable_enable_r = main_genericstandalone_interface1_csr_bus_dat_w[0];
assign main_genericstandalone_dma_enable_enable_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 1'd0));
assign main_genericstandalone_base_address1_r = main_genericstandalone_interface1_csr_bus_dat_w[0];
assign main_genericstandalone_base_address1_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 1'd1));
assign main_genericstandalone_base_address0_r = main_genericstandalone_interface1_csr_bus_dat_w[31:0];
assign main_genericstandalone_base_address0_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 2'd2));
assign main_genericstandalone_time_offset1_r = main_genericstandalone_interface1_csr_bus_dat_w[31:0];
assign main_genericstandalone_time_offset1_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 2'd3));
assign main_genericstandalone_time_offset0_r = main_genericstandalone_interface1_csr_bus_dat_w[31:0];
assign main_genericstandalone_time_offset0_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 3'd4));
assign main_genericstandalone_dma_cri_master_error_r = main_genericstandalone_interface1_csr_bus_dat_w[1:0];
assign main_genericstandalone_dma_cri_master_error_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 3'd5));
assign main_genericstandalone_error_channel_r = main_genericstandalone_interface1_csr_bus_dat_w[23:0];
assign main_genericstandalone_error_channel_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 3'd6));
assign main_genericstandalone_error_timestamp1_r = main_genericstandalone_interface1_csr_bus_dat_w[31:0];
assign main_genericstandalone_error_timestamp1_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 3'd7));
assign main_genericstandalone_error_timestamp0_r = main_genericstandalone_interface1_csr_bus_dat_w[31:0];
assign main_genericstandalone_error_timestamp0_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 4'd8));
assign main_genericstandalone_error_address_r = main_genericstandalone_interface1_csr_bus_dat_w[15:0];
assign main_genericstandalone_error_address_re = ((((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb) & (~main_genericstandalone_interface1_csr_bus_ack)) & main_genericstandalone_interface1_csr_bus_we) & (main_genericstandalone_interface1_csr_bus_adr[3:0] == 4'd9));
assign main_genericstandalone_dma_dma_storage = main_genericstandalone_dma_dma_storage_full[32:4];
assign main_genericstandalone_base_address1_w = main_genericstandalone_dma_dma_storage_full[32];
assign main_genericstandalone_base_address0_w = {main_genericstandalone_dma_dma_storage_full[31:4], {28{1'd0}}};
assign main_genericstandalone_dma_time_offset_storage = main_genericstandalone_dma_time_offset_storage_full[63:0];
assign main_genericstandalone_time_offset1_w = main_genericstandalone_dma_time_offset_storage_full[63:32];
assign main_genericstandalone_time_offset0_w = main_genericstandalone_dma_time_offset_storage_full[31:0];
assign main_genericstandalone_error_channel_w = main_genericstandalone_dma_cri_master_error_channel_status[23:0];
assign main_genericstandalone_error_timestamp1_w = main_genericstandalone_dma_cri_master_error_timestamp_status[63:32];
assign main_genericstandalone_error_timestamp0_w = main_genericstandalone_dma_cri_master_error_timestamp_status[31:0];
assign main_genericstandalone_error_address_w = main_genericstandalone_dma_cri_master_error_address_status[15:0];
assign main_genericstandalone_cri_con_shared_cmd = builder_comb_rhs_self11;
assign main_genericstandalone_cri_con_shared_chan_sel = builder_comb_rhs_self12;
assign main_genericstandalone_cri_con_shared_o_timestamp = builder_comb_rhs_self13;
assign main_genericstandalone_cri_con_shared_o_data = builder_comb_rhs_self14;
assign main_genericstandalone_cri_con_shared_o_address = builder_comb_rhs_self15;
assign main_genericstandalone_cri_con_shared_i_timeout = builder_comb_rhs_self16;
assign main_genericstandalone_rtio_cri_o_status = main_genericstandalone_cri_con_shared_o_status;
assign main_genericstandalone_dma_cri_master_cri_o_status = main_genericstandalone_cri_con_shared_o_status;
assign main_genericstandalone_rtio_cri_o_buffer_space_valid = main_genericstandalone_cri_con_shared_o_buffer_space_valid;
assign main_genericstandalone_dma_cri_master_cri_o_buffer_space_valid = main_genericstandalone_cri_con_shared_o_buffer_space_valid;
assign main_genericstandalone_rtio_cri_o_buffer_space = main_genericstandalone_cri_con_shared_o_buffer_space;
assign main_genericstandalone_dma_cri_master_cri_o_buffer_space = main_genericstandalone_cri_con_shared_o_buffer_space;
assign main_genericstandalone_rtio_cri_i_data = main_genericstandalone_cri_con_shared_i_data;
assign main_genericstandalone_dma_cri_master_cri_i_data = main_genericstandalone_cri_con_shared_i_data;
assign main_genericstandalone_rtio_cri_i_timestamp = main_genericstandalone_cri_con_shared_i_timestamp;
assign main_genericstandalone_dma_cri_master_cri_i_timestamp = main_genericstandalone_cri_con_shared_i_timestamp;
assign main_genericstandalone_rtio_cri_i_status = main_genericstandalone_cri_con_shared_i_status;
assign main_genericstandalone_dma_cri_master_cri_i_status = main_genericstandalone_cri_con_shared_i_status;
assign main_genericstandalone_rtio_core_cri_chan_sel = main_genericstandalone_cri_con_shared_chan_sel;
assign main_genericstandalone_rtio_core_cri_o_timestamp = main_genericstandalone_cri_con_shared_o_timestamp;
assign main_genericstandalone_rtio_core_cri_o_data = main_genericstandalone_cri_con_shared_o_data;
assign main_genericstandalone_rtio_core_cri_o_address = main_genericstandalone_cri_con_shared_o_address;
assign main_genericstandalone_rtio_core_cri_i_timeout = main_genericstandalone_cri_con_shared_i_timeout;

// synthesis translate_off
reg dummy_d_210;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_core_cri_cmd <= 2'd0;
	if ((main_genericstandalone_cri_con_selected == 1'd0)) begin
		main_genericstandalone_rtio_core_cri_cmd <= main_genericstandalone_cri_con_shared_cmd;
	end
// synthesis translate_off
	dummy_d_210 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_211;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_cri_con_shared_o_status <= 3'd0;
	main_genericstandalone_cri_con_shared_o_buffer_space_valid <= 1'd0;
	main_genericstandalone_cri_con_shared_o_buffer_space <= 16'd0;
	main_genericstandalone_cri_con_shared_i_data <= 32'd0;
	main_genericstandalone_cri_con_shared_i_timestamp <= 64'd0;
	main_genericstandalone_cri_con_shared_i_status <= 4'd0;
	case (main_genericstandalone_cri_con_selected)
		1'd0: begin
			main_genericstandalone_cri_con_shared_o_status <= main_genericstandalone_rtio_core_cri_o_status;
			main_genericstandalone_cri_con_shared_o_buffer_space_valid <= main_genericstandalone_rtio_core_cri_o_buffer_space_valid;
			main_genericstandalone_cri_con_shared_o_buffer_space <= main_genericstandalone_rtio_core_cri_o_buffer_space;
			main_genericstandalone_cri_con_shared_i_data <= main_genericstandalone_rtio_core_cri_i_data;
			main_genericstandalone_cri_con_shared_i_timestamp <= main_genericstandalone_rtio_core_cri_i_timestamp;
			main_genericstandalone_cri_con_shared_i_status <= main_genericstandalone_rtio_core_cri_i_status;
		end
	endcase
// synthesis translate_off
	dummy_d_211 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_selected0_r = main_genericstandalone_interface2_csr_bus_dat_w[1:0];
assign main_genericstandalone_selected0_re = ((((main_genericstandalone_interface2_csr_bus_cyc & main_genericstandalone_interface2_csr_bus_stb) & (~main_genericstandalone_interface2_csr_bus_ack)) & main_genericstandalone_interface2_csr_bus_we) & (main_genericstandalone_interface2_csr_bus_adr[0] == 1'd0));
assign main_genericstandalone_cri_con_storage = main_genericstandalone_cri_con_storage_full[1:0];
assign main_genericstandalone_selected0_w = main_genericstandalone_cri_con_storage_full[1:0];
assign main_genericstandalone_mon_bussynchronizer0_i = main_inout_8x0_serdes_i0[7];
assign main_genericstandalone_mon_bussynchronizer1_i = main_inout_8x0_serdes_oe;
assign main_genericstandalone_mon_bussynchronizer2_i = main_inout_8x1_serdes_i0[7];
assign main_genericstandalone_mon_bussynchronizer3_i = main_inout_8x1_serdes_oe;
assign main_genericstandalone_mon_bussynchronizer4_i = main_inout_8x2_serdes_i0[7];
assign main_genericstandalone_mon_bussynchronizer5_i = main_inout_8x2_serdes_oe;
assign main_genericstandalone_mon_bussynchronizer6_i = main_inout_8x3_serdes_i0[7];
assign main_genericstandalone_mon_bussynchronizer7_i = main_inout_8x3_serdes_oe;
assign main_genericstandalone_mon_bussynchronizer8_i = main_output_8x0_o0[7];
assign main_genericstandalone_mon_bussynchronizer9_i = main_output_8x1_o0[7];
assign main_genericstandalone_mon_bussynchronizer10_i = main_output_8x2_o[7];
assign main_genericstandalone_mon_bussynchronizer11_i = main_output_8x3_o[7];
assign main_genericstandalone_mon_bussynchronizer12_i = main_output_8x4_o[7];
assign main_genericstandalone_mon_bussynchronizer13_i = main_output_8x5_o[7];
assign main_genericstandalone_mon_bussynchronizer14_i = main_output_8x6_o[7];
assign main_genericstandalone_mon_bussynchronizer15_i = main_output_8x7_o[7];
assign main_genericstandalone_mon_bussynchronizer16_i = main_output_8x8_o[7];
assign main_genericstandalone_mon_bussynchronizer17_i = main_output_8x9_o[7];
assign main_genericstandalone_mon_bussynchronizer18_i = main_output_8x10_o[7];
assign main_genericstandalone_mon_bussynchronizer19_i = main_output_8x11_o[7];
assign main_genericstandalone_mon_bussynchronizer20_i = main_urukulmonitor00;
assign main_genericstandalone_mon_bussynchronizer21_i = main_urukulmonitor01;
assign main_genericstandalone_mon_bussynchronizer22_i = main_urukulmonitor02;
assign main_genericstandalone_mon_bussynchronizer23_i = main_urukulmonitor03;
assign main_genericstandalone_mon_bussynchronizer24_i = main_output_8x0_o1[7];
assign main_genericstandalone_mon_bussynchronizer25_i = main_output_8x12_o[7];
assign main_genericstandalone_mon_bussynchronizer26_i = main_output_8x13_o[7];
assign main_genericstandalone_mon_bussynchronizer27_i = main_output_8x14_o[7];
assign main_genericstandalone_mon_bussynchronizer28_i = main_output_8x15_o[7];
assign main_genericstandalone_mon_bussynchronizer29_i = main_urukulmonitor10;
assign main_genericstandalone_mon_bussynchronizer30_i = main_urukulmonitor11;
assign main_genericstandalone_mon_bussynchronizer31_i = main_urukulmonitor12;
assign main_genericstandalone_mon_bussynchronizer32_i = main_urukulmonitor13;
assign main_genericstandalone_mon_bussynchronizer33_i = main_output_8x1_o1[7];
assign main_genericstandalone_mon_bussynchronizer34_i = main_output_8x16_o[7];
assign main_genericstandalone_mon_bussynchronizer35_i = main_output_8x17_o[7];
assign main_genericstandalone_mon_bussynchronizer36_i = main_output_8x18_o[7];
assign main_genericstandalone_mon_bussynchronizer37_i = main_output_8x19_o[7];
assign main_genericstandalone_mon_bussynchronizer38_i = main_output_8x20_o[7];
assign main_genericstandalone_mon_bussynchronizer39_i = main_ad53xxmonitor0;
assign main_genericstandalone_mon_bussynchronizer40_i = main_ad53xxmonitor1;
assign main_genericstandalone_mon_bussynchronizer41_i = main_ad53xxmonitor2;
assign main_genericstandalone_mon_bussynchronizer42_i = main_ad53xxmonitor3;
assign main_genericstandalone_mon_bussynchronizer43_i = main_ad53xxmonitor4;
assign main_genericstandalone_mon_bussynchronizer44_i = main_ad53xxmonitor5;
assign main_genericstandalone_mon_bussynchronizer45_i = main_ad53xxmonitor6;
assign main_genericstandalone_mon_bussynchronizer46_i = main_ad53xxmonitor7;
assign main_genericstandalone_mon_bussynchronizer47_i = main_ad53xxmonitor8;
assign main_genericstandalone_mon_bussynchronizer48_i = main_ad53xxmonitor9;
assign main_genericstandalone_mon_bussynchronizer49_i = main_ad53xxmonitor10;
assign main_genericstandalone_mon_bussynchronizer50_i = main_ad53xxmonitor11;
assign main_genericstandalone_mon_bussynchronizer51_i = main_ad53xxmonitor12;
assign main_genericstandalone_mon_bussynchronizer52_i = main_ad53xxmonitor13;
assign main_genericstandalone_mon_bussynchronizer53_i = main_ad53xxmonitor14;
assign main_genericstandalone_mon_bussynchronizer54_i = main_ad53xxmonitor15;
assign main_genericstandalone_mon_bussynchronizer55_i = main_ad53xxmonitor16;
assign main_genericstandalone_mon_bussynchronizer56_i = main_ad53xxmonitor17;
assign main_genericstandalone_mon_bussynchronizer57_i = main_ad53xxmonitor18;
assign main_genericstandalone_mon_bussynchronizer58_i = main_ad53xxmonitor19;
assign main_genericstandalone_mon_bussynchronizer59_i = main_ad53xxmonitor20;
assign main_genericstandalone_mon_bussynchronizer60_i = main_ad53xxmonitor21;
assign main_genericstandalone_mon_bussynchronizer61_i = main_ad53xxmonitor22;
assign main_genericstandalone_mon_bussynchronizer62_i = main_ad53xxmonitor23;
assign main_genericstandalone_mon_bussynchronizer63_i = main_ad53xxmonitor24;
assign main_genericstandalone_mon_bussynchronizer64_i = main_ad53xxmonitor25;
assign main_genericstandalone_mon_bussynchronizer65_i = main_ad53xxmonitor26;
assign main_genericstandalone_mon_bussynchronizer66_i = main_ad53xxmonitor27;
assign main_genericstandalone_mon_bussynchronizer67_i = main_ad53xxmonitor28;
assign main_genericstandalone_mon_bussynchronizer68_i = main_ad53xxmonitor29;
assign main_genericstandalone_mon_bussynchronizer69_i = main_ad53xxmonitor30;
assign main_genericstandalone_mon_bussynchronizer70_i = main_ad53xxmonitor31;
assign main_genericstandalone_mon_bussynchronizer71_i = main_ldac_phy_o[7];
assign main_genericstandalone_mon_bussynchronizer72_i = main_clr_phy_o[7];
assign main_genericstandalone_mon_bussynchronizer73_i = main_output0_pad_o;
assign main_genericstandalone_mon_bussynchronizer74_i = main_output1_pad_o;
assign main_genericstandalone_mon_bussynchronizer75_i = main_output2_pad_o;
assign main_genericstandalone_mon_bussynchronizer20_wait = (~main_genericstandalone_mon_bussynchronizer20_ping_i);
assign main_genericstandalone_mon_bussynchronizer20_ping_i = ((main_genericstandalone_mon_bussynchronizer20_starter | main_genericstandalone_mon_bussynchronizer20_pong_o) | main_genericstandalone_mon_bussynchronizer20_done);
assign main_genericstandalone_mon_bussynchronizer20_pong_i = main_genericstandalone_mon_bussynchronizer20_ping_o1;
assign main_genericstandalone_mon_bussynchronizer20_ping_o0 = (main_genericstandalone_mon_bussynchronizer20_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer20_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer20_pong_o = (main_genericstandalone_mon_bussynchronizer20_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer20_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer20_done = (main_genericstandalone_mon_bussynchronizer20_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer21_wait = (~main_genericstandalone_mon_bussynchronizer21_ping_i);
assign main_genericstandalone_mon_bussynchronizer21_ping_i = ((main_genericstandalone_mon_bussynchronizer21_starter | main_genericstandalone_mon_bussynchronizer21_pong_o) | main_genericstandalone_mon_bussynchronizer21_done);
assign main_genericstandalone_mon_bussynchronizer21_pong_i = main_genericstandalone_mon_bussynchronizer21_ping_o1;
assign main_genericstandalone_mon_bussynchronizer21_ping_o0 = (main_genericstandalone_mon_bussynchronizer21_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer21_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer21_pong_o = (main_genericstandalone_mon_bussynchronizer21_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer21_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer21_done = (main_genericstandalone_mon_bussynchronizer21_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer22_wait = (~main_genericstandalone_mon_bussynchronizer22_ping_i);
assign main_genericstandalone_mon_bussynchronizer22_ping_i = ((main_genericstandalone_mon_bussynchronizer22_starter | main_genericstandalone_mon_bussynchronizer22_pong_o) | main_genericstandalone_mon_bussynchronizer22_done);
assign main_genericstandalone_mon_bussynchronizer22_pong_i = main_genericstandalone_mon_bussynchronizer22_ping_o1;
assign main_genericstandalone_mon_bussynchronizer22_ping_o0 = (main_genericstandalone_mon_bussynchronizer22_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer22_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer22_pong_o = (main_genericstandalone_mon_bussynchronizer22_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer22_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer22_done = (main_genericstandalone_mon_bussynchronizer22_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer23_wait = (~main_genericstandalone_mon_bussynchronizer23_ping_i);
assign main_genericstandalone_mon_bussynchronizer23_ping_i = ((main_genericstandalone_mon_bussynchronizer23_starter | main_genericstandalone_mon_bussynchronizer23_pong_o) | main_genericstandalone_mon_bussynchronizer23_done);
assign main_genericstandalone_mon_bussynchronizer23_pong_i = main_genericstandalone_mon_bussynchronizer23_ping_o1;
assign main_genericstandalone_mon_bussynchronizer23_ping_o0 = (main_genericstandalone_mon_bussynchronizer23_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer23_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer23_pong_o = (main_genericstandalone_mon_bussynchronizer23_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer23_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer23_done = (main_genericstandalone_mon_bussynchronizer23_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer29_wait = (~main_genericstandalone_mon_bussynchronizer29_ping_i);
assign main_genericstandalone_mon_bussynchronizer29_ping_i = ((main_genericstandalone_mon_bussynchronizer29_starter | main_genericstandalone_mon_bussynchronizer29_pong_o) | main_genericstandalone_mon_bussynchronizer29_done);
assign main_genericstandalone_mon_bussynchronizer29_pong_i = main_genericstandalone_mon_bussynchronizer29_ping_o1;
assign main_genericstandalone_mon_bussynchronizer29_ping_o0 = (main_genericstandalone_mon_bussynchronizer29_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer29_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer29_pong_o = (main_genericstandalone_mon_bussynchronizer29_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer29_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer29_done = (main_genericstandalone_mon_bussynchronizer29_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer30_wait = (~main_genericstandalone_mon_bussynchronizer30_ping_i);
assign main_genericstandalone_mon_bussynchronizer30_ping_i = ((main_genericstandalone_mon_bussynchronizer30_starter | main_genericstandalone_mon_bussynchronizer30_pong_o) | main_genericstandalone_mon_bussynchronizer30_done);
assign main_genericstandalone_mon_bussynchronizer30_pong_i = main_genericstandalone_mon_bussynchronizer30_ping_o1;
assign main_genericstandalone_mon_bussynchronizer30_ping_o0 = (main_genericstandalone_mon_bussynchronizer30_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer30_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer30_pong_o = (main_genericstandalone_mon_bussynchronizer30_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer30_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer30_done = (main_genericstandalone_mon_bussynchronizer30_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer31_wait = (~main_genericstandalone_mon_bussynchronizer31_ping_i);
assign main_genericstandalone_mon_bussynchronizer31_ping_i = ((main_genericstandalone_mon_bussynchronizer31_starter | main_genericstandalone_mon_bussynchronizer31_pong_o) | main_genericstandalone_mon_bussynchronizer31_done);
assign main_genericstandalone_mon_bussynchronizer31_pong_i = main_genericstandalone_mon_bussynchronizer31_ping_o1;
assign main_genericstandalone_mon_bussynchronizer31_ping_o0 = (main_genericstandalone_mon_bussynchronizer31_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer31_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer31_pong_o = (main_genericstandalone_mon_bussynchronizer31_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer31_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer31_done = (main_genericstandalone_mon_bussynchronizer31_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer32_wait = (~main_genericstandalone_mon_bussynchronizer32_ping_i);
assign main_genericstandalone_mon_bussynchronizer32_ping_i = ((main_genericstandalone_mon_bussynchronizer32_starter | main_genericstandalone_mon_bussynchronizer32_pong_o) | main_genericstandalone_mon_bussynchronizer32_done);
assign main_genericstandalone_mon_bussynchronizer32_pong_i = main_genericstandalone_mon_bussynchronizer32_ping_o1;
assign main_genericstandalone_mon_bussynchronizer32_ping_o0 = (main_genericstandalone_mon_bussynchronizer32_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer32_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer32_pong_o = (main_genericstandalone_mon_bussynchronizer32_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer32_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer32_done = (main_genericstandalone_mon_bussynchronizer32_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer39_wait = (~main_genericstandalone_mon_bussynchronizer39_ping_i);
assign main_genericstandalone_mon_bussynchronizer39_ping_i = ((main_genericstandalone_mon_bussynchronizer39_starter | main_genericstandalone_mon_bussynchronizer39_pong_o) | main_genericstandalone_mon_bussynchronizer39_done);
assign main_genericstandalone_mon_bussynchronizer39_pong_i = main_genericstandalone_mon_bussynchronizer39_ping_o1;
assign main_genericstandalone_mon_bussynchronizer39_ping_o0 = (main_genericstandalone_mon_bussynchronizer39_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer39_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer39_pong_o = (main_genericstandalone_mon_bussynchronizer39_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer39_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer39_done = (main_genericstandalone_mon_bussynchronizer39_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer40_wait = (~main_genericstandalone_mon_bussynchronizer40_ping_i);
assign main_genericstandalone_mon_bussynchronizer40_ping_i = ((main_genericstandalone_mon_bussynchronizer40_starter | main_genericstandalone_mon_bussynchronizer40_pong_o) | main_genericstandalone_mon_bussynchronizer40_done);
assign main_genericstandalone_mon_bussynchronizer40_pong_i = main_genericstandalone_mon_bussynchronizer40_ping_o1;
assign main_genericstandalone_mon_bussynchronizer40_ping_o0 = (main_genericstandalone_mon_bussynchronizer40_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer40_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer40_pong_o = (main_genericstandalone_mon_bussynchronizer40_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer40_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer40_done = (main_genericstandalone_mon_bussynchronizer40_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer41_wait = (~main_genericstandalone_mon_bussynchronizer41_ping_i);
assign main_genericstandalone_mon_bussynchronizer41_ping_i = ((main_genericstandalone_mon_bussynchronizer41_starter | main_genericstandalone_mon_bussynchronizer41_pong_o) | main_genericstandalone_mon_bussynchronizer41_done);
assign main_genericstandalone_mon_bussynchronizer41_pong_i = main_genericstandalone_mon_bussynchronizer41_ping_o1;
assign main_genericstandalone_mon_bussynchronizer41_ping_o0 = (main_genericstandalone_mon_bussynchronizer41_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer41_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer41_pong_o = (main_genericstandalone_mon_bussynchronizer41_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer41_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer41_done = (main_genericstandalone_mon_bussynchronizer41_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer42_wait = (~main_genericstandalone_mon_bussynchronizer42_ping_i);
assign main_genericstandalone_mon_bussynchronizer42_ping_i = ((main_genericstandalone_mon_bussynchronizer42_starter | main_genericstandalone_mon_bussynchronizer42_pong_o) | main_genericstandalone_mon_bussynchronizer42_done);
assign main_genericstandalone_mon_bussynchronizer42_pong_i = main_genericstandalone_mon_bussynchronizer42_ping_o1;
assign main_genericstandalone_mon_bussynchronizer42_ping_o0 = (main_genericstandalone_mon_bussynchronizer42_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer42_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer42_pong_o = (main_genericstandalone_mon_bussynchronizer42_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer42_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer42_done = (main_genericstandalone_mon_bussynchronizer42_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer43_wait = (~main_genericstandalone_mon_bussynchronizer43_ping_i);
assign main_genericstandalone_mon_bussynchronizer43_ping_i = ((main_genericstandalone_mon_bussynchronizer43_starter | main_genericstandalone_mon_bussynchronizer43_pong_o) | main_genericstandalone_mon_bussynchronizer43_done);
assign main_genericstandalone_mon_bussynchronizer43_pong_i = main_genericstandalone_mon_bussynchronizer43_ping_o1;
assign main_genericstandalone_mon_bussynchronizer43_ping_o0 = (main_genericstandalone_mon_bussynchronizer43_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer43_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer43_pong_o = (main_genericstandalone_mon_bussynchronizer43_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer43_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer43_done = (main_genericstandalone_mon_bussynchronizer43_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer44_wait = (~main_genericstandalone_mon_bussynchronizer44_ping_i);
assign main_genericstandalone_mon_bussynchronizer44_ping_i = ((main_genericstandalone_mon_bussynchronizer44_starter | main_genericstandalone_mon_bussynchronizer44_pong_o) | main_genericstandalone_mon_bussynchronizer44_done);
assign main_genericstandalone_mon_bussynchronizer44_pong_i = main_genericstandalone_mon_bussynchronizer44_ping_o1;
assign main_genericstandalone_mon_bussynchronizer44_ping_o0 = (main_genericstandalone_mon_bussynchronizer44_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer44_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer44_pong_o = (main_genericstandalone_mon_bussynchronizer44_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer44_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer44_done = (main_genericstandalone_mon_bussynchronizer44_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer45_wait = (~main_genericstandalone_mon_bussynchronizer45_ping_i);
assign main_genericstandalone_mon_bussynchronizer45_ping_i = ((main_genericstandalone_mon_bussynchronizer45_starter | main_genericstandalone_mon_bussynchronizer45_pong_o) | main_genericstandalone_mon_bussynchronizer45_done);
assign main_genericstandalone_mon_bussynchronizer45_pong_i = main_genericstandalone_mon_bussynchronizer45_ping_o1;
assign main_genericstandalone_mon_bussynchronizer45_ping_o0 = (main_genericstandalone_mon_bussynchronizer45_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer45_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer45_pong_o = (main_genericstandalone_mon_bussynchronizer45_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer45_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer45_done = (main_genericstandalone_mon_bussynchronizer45_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer46_wait = (~main_genericstandalone_mon_bussynchronizer46_ping_i);
assign main_genericstandalone_mon_bussynchronizer46_ping_i = ((main_genericstandalone_mon_bussynchronizer46_starter | main_genericstandalone_mon_bussynchronizer46_pong_o) | main_genericstandalone_mon_bussynchronizer46_done);
assign main_genericstandalone_mon_bussynchronizer46_pong_i = main_genericstandalone_mon_bussynchronizer46_ping_o1;
assign main_genericstandalone_mon_bussynchronizer46_ping_o0 = (main_genericstandalone_mon_bussynchronizer46_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer46_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer46_pong_o = (main_genericstandalone_mon_bussynchronizer46_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer46_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer46_done = (main_genericstandalone_mon_bussynchronizer46_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer47_wait = (~main_genericstandalone_mon_bussynchronizer47_ping_i);
assign main_genericstandalone_mon_bussynchronizer47_ping_i = ((main_genericstandalone_mon_bussynchronizer47_starter | main_genericstandalone_mon_bussynchronizer47_pong_o) | main_genericstandalone_mon_bussynchronizer47_done);
assign main_genericstandalone_mon_bussynchronizer47_pong_i = main_genericstandalone_mon_bussynchronizer47_ping_o1;
assign main_genericstandalone_mon_bussynchronizer47_ping_o0 = (main_genericstandalone_mon_bussynchronizer47_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer47_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer47_pong_o = (main_genericstandalone_mon_bussynchronizer47_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer47_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer47_done = (main_genericstandalone_mon_bussynchronizer47_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer48_wait = (~main_genericstandalone_mon_bussynchronizer48_ping_i);
assign main_genericstandalone_mon_bussynchronizer48_ping_i = ((main_genericstandalone_mon_bussynchronizer48_starter | main_genericstandalone_mon_bussynchronizer48_pong_o) | main_genericstandalone_mon_bussynchronizer48_done);
assign main_genericstandalone_mon_bussynchronizer48_pong_i = main_genericstandalone_mon_bussynchronizer48_ping_o1;
assign main_genericstandalone_mon_bussynchronizer48_ping_o0 = (main_genericstandalone_mon_bussynchronizer48_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer48_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer48_pong_o = (main_genericstandalone_mon_bussynchronizer48_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer48_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer48_done = (main_genericstandalone_mon_bussynchronizer48_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer49_wait = (~main_genericstandalone_mon_bussynchronizer49_ping_i);
assign main_genericstandalone_mon_bussynchronizer49_ping_i = ((main_genericstandalone_mon_bussynchronizer49_starter | main_genericstandalone_mon_bussynchronizer49_pong_o) | main_genericstandalone_mon_bussynchronizer49_done);
assign main_genericstandalone_mon_bussynchronizer49_pong_i = main_genericstandalone_mon_bussynchronizer49_ping_o1;
assign main_genericstandalone_mon_bussynchronizer49_ping_o0 = (main_genericstandalone_mon_bussynchronizer49_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer49_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer49_pong_o = (main_genericstandalone_mon_bussynchronizer49_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer49_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer49_done = (main_genericstandalone_mon_bussynchronizer49_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer50_wait = (~main_genericstandalone_mon_bussynchronizer50_ping_i);
assign main_genericstandalone_mon_bussynchronizer50_ping_i = ((main_genericstandalone_mon_bussynchronizer50_starter | main_genericstandalone_mon_bussynchronizer50_pong_o) | main_genericstandalone_mon_bussynchronizer50_done);
assign main_genericstandalone_mon_bussynchronizer50_pong_i = main_genericstandalone_mon_bussynchronizer50_ping_o1;
assign main_genericstandalone_mon_bussynchronizer50_ping_o0 = (main_genericstandalone_mon_bussynchronizer50_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer50_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer50_pong_o = (main_genericstandalone_mon_bussynchronizer50_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer50_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer50_done = (main_genericstandalone_mon_bussynchronizer50_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer51_wait = (~main_genericstandalone_mon_bussynchronizer51_ping_i);
assign main_genericstandalone_mon_bussynchronizer51_ping_i = ((main_genericstandalone_mon_bussynchronizer51_starter | main_genericstandalone_mon_bussynchronizer51_pong_o) | main_genericstandalone_mon_bussynchronizer51_done);
assign main_genericstandalone_mon_bussynchronizer51_pong_i = main_genericstandalone_mon_bussynchronizer51_ping_o1;
assign main_genericstandalone_mon_bussynchronizer51_ping_o0 = (main_genericstandalone_mon_bussynchronizer51_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer51_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer51_pong_o = (main_genericstandalone_mon_bussynchronizer51_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer51_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer51_done = (main_genericstandalone_mon_bussynchronizer51_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer52_wait = (~main_genericstandalone_mon_bussynchronizer52_ping_i);
assign main_genericstandalone_mon_bussynchronizer52_ping_i = ((main_genericstandalone_mon_bussynchronizer52_starter | main_genericstandalone_mon_bussynchronizer52_pong_o) | main_genericstandalone_mon_bussynchronizer52_done);
assign main_genericstandalone_mon_bussynchronizer52_pong_i = main_genericstandalone_mon_bussynchronizer52_ping_o1;
assign main_genericstandalone_mon_bussynchronizer52_ping_o0 = (main_genericstandalone_mon_bussynchronizer52_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer52_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer52_pong_o = (main_genericstandalone_mon_bussynchronizer52_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer52_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer52_done = (main_genericstandalone_mon_bussynchronizer52_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer53_wait = (~main_genericstandalone_mon_bussynchronizer53_ping_i);
assign main_genericstandalone_mon_bussynchronizer53_ping_i = ((main_genericstandalone_mon_bussynchronizer53_starter | main_genericstandalone_mon_bussynchronizer53_pong_o) | main_genericstandalone_mon_bussynchronizer53_done);
assign main_genericstandalone_mon_bussynchronizer53_pong_i = main_genericstandalone_mon_bussynchronizer53_ping_o1;
assign main_genericstandalone_mon_bussynchronizer53_ping_o0 = (main_genericstandalone_mon_bussynchronizer53_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer53_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer53_pong_o = (main_genericstandalone_mon_bussynchronizer53_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer53_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer53_done = (main_genericstandalone_mon_bussynchronizer53_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer54_wait = (~main_genericstandalone_mon_bussynchronizer54_ping_i);
assign main_genericstandalone_mon_bussynchronizer54_ping_i = ((main_genericstandalone_mon_bussynchronizer54_starter | main_genericstandalone_mon_bussynchronizer54_pong_o) | main_genericstandalone_mon_bussynchronizer54_done);
assign main_genericstandalone_mon_bussynchronizer54_pong_i = main_genericstandalone_mon_bussynchronizer54_ping_o1;
assign main_genericstandalone_mon_bussynchronizer54_ping_o0 = (main_genericstandalone_mon_bussynchronizer54_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer54_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer54_pong_o = (main_genericstandalone_mon_bussynchronizer54_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer54_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer54_done = (main_genericstandalone_mon_bussynchronizer54_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer55_wait = (~main_genericstandalone_mon_bussynchronizer55_ping_i);
assign main_genericstandalone_mon_bussynchronizer55_ping_i = ((main_genericstandalone_mon_bussynchronizer55_starter | main_genericstandalone_mon_bussynchronizer55_pong_o) | main_genericstandalone_mon_bussynchronizer55_done);
assign main_genericstandalone_mon_bussynchronizer55_pong_i = main_genericstandalone_mon_bussynchronizer55_ping_o1;
assign main_genericstandalone_mon_bussynchronizer55_ping_o0 = (main_genericstandalone_mon_bussynchronizer55_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer55_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer55_pong_o = (main_genericstandalone_mon_bussynchronizer55_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer55_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer55_done = (main_genericstandalone_mon_bussynchronizer55_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer56_wait = (~main_genericstandalone_mon_bussynchronizer56_ping_i);
assign main_genericstandalone_mon_bussynchronizer56_ping_i = ((main_genericstandalone_mon_bussynchronizer56_starter | main_genericstandalone_mon_bussynchronizer56_pong_o) | main_genericstandalone_mon_bussynchronizer56_done);
assign main_genericstandalone_mon_bussynchronizer56_pong_i = main_genericstandalone_mon_bussynchronizer56_ping_o1;
assign main_genericstandalone_mon_bussynchronizer56_ping_o0 = (main_genericstandalone_mon_bussynchronizer56_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer56_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer56_pong_o = (main_genericstandalone_mon_bussynchronizer56_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer56_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer56_done = (main_genericstandalone_mon_bussynchronizer56_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer57_wait = (~main_genericstandalone_mon_bussynchronizer57_ping_i);
assign main_genericstandalone_mon_bussynchronizer57_ping_i = ((main_genericstandalone_mon_bussynchronizer57_starter | main_genericstandalone_mon_bussynchronizer57_pong_o) | main_genericstandalone_mon_bussynchronizer57_done);
assign main_genericstandalone_mon_bussynchronizer57_pong_i = main_genericstandalone_mon_bussynchronizer57_ping_o1;
assign main_genericstandalone_mon_bussynchronizer57_ping_o0 = (main_genericstandalone_mon_bussynchronizer57_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer57_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer57_pong_o = (main_genericstandalone_mon_bussynchronizer57_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer57_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer57_done = (main_genericstandalone_mon_bussynchronizer57_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer58_wait = (~main_genericstandalone_mon_bussynchronizer58_ping_i);
assign main_genericstandalone_mon_bussynchronizer58_ping_i = ((main_genericstandalone_mon_bussynchronizer58_starter | main_genericstandalone_mon_bussynchronizer58_pong_o) | main_genericstandalone_mon_bussynchronizer58_done);
assign main_genericstandalone_mon_bussynchronizer58_pong_i = main_genericstandalone_mon_bussynchronizer58_ping_o1;
assign main_genericstandalone_mon_bussynchronizer58_ping_o0 = (main_genericstandalone_mon_bussynchronizer58_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer58_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer58_pong_o = (main_genericstandalone_mon_bussynchronizer58_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer58_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer58_done = (main_genericstandalone_mon_bussynchronizer58_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer59_wait = (~main_genericstandalone_mon_bussynchronizer59_ping_i);
assign main_genericstandalone_mon_bussynchronizer59_ping_i = ((main_genericstandalone_mon_bussynchronizer59_starter | main_genericstandalone_mon_bussynchronizer59_pong_o) | main_genericstandalone_mon_bussynchronizer59_done);
assign main_genericstandalone_mon_bussynchronizer59_pong_i = main_genericstandalone_mon_bussynchronizer59_ping_o1;
assign main_genericstandalone_mon_bussynchronizer59_ping_o0 = (main_genericstandalone_mon_bussynchronizer59_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer59_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer59_pong_o = (main_genericstandalone_mon_bussynchronizer59_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer59_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer59_done = (main_genericstandalone_mon_bussynchronizer59_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer60_wait = (~main_genericstandalone_mon_bussynchronizer60_ping_i);
assign main_genericstandalone_mon_bussynchronizer60_ping_i = ((main_genericstandalone_mon_bussynchronizer60_starter | main_genericstandalone_mon_bussynchronizer60_pong_o) | main_genericstandalone_mon_bussynchronizer60_done);
assign main_genericstandalone_mon_bussynchronizer60_pong_i = main_genericstandalone_mon_bussynchronizer60_ping_o1;
assign main_genericstandalone_mon_bussynchronizer60_ping_o0 = (main_genericstandalone_mon_bussynchronizer60_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer60_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer60_pong_o = (main_genericstandalone_mon_bussynchronizer60_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer60_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer60_done = (main_genericstandalone_mon_bussynchronizer60_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer61_wait = (~main_genericstandalone_mon_bussynchronizer61_ping_i);
assign main_genericstandalone_mon_bussynchronizer61_ping_i = ((main_genericstandalone_mon_bussynchronizer61_starter | main_genericstandalone_mon_bussynchronizer61_pong_o) | main_genericstandalone_mon_bussynchronizer61_done);
assign main_genericstandalone_mon_bussynchronizer61_pong_i = main_genericstandalone_mon_bussynchronizer61_ping_o1;
assign main_genericstandalone_mon_bussynchronizer61_ping_o0 = (main_genericstandalone_mon_bussynchronizer61_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer61_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer61_pong_o = (main_genericstandalone_mon_bussynchronizer61_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer61_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer61_done = (main_genericstandalone_mon_bussynchronizer61_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer62_wait = (~main_genericstandalone_mon_bussynchronizer62_ping_i);
assign main_genericstandalone_mon_bussynchronizer62_ping_i = ((main_genericstandalone_mon_bussynchronizer62_starter | main_genericstandalone_mon_bussynchronizer62_pong_o) | main_genericstandalone_mon_bussynchronizer62_done);
assign main_genericstandalone_mon_bussynchronizer62_pong_i = main_genericstandalone_mon_bussynchronizer62_ping_o1;
assign main_genericstandalone_mon_bussynchronizer62_ping_o0 = (main_genericstandalone_mon_bussynchronizer62_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer62_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer62_pong_o = (main_genericstandalone_mon_bussynchronizer62_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer62_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer62_done = (main_genericstandalone_mon_bussynchronizer62_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer63_wait = (~main_genericstandalone_mon_bussynchronizer63_ping_i);
assign main_genericstandalone_mon_bussynchronizer63_ping_i = ((main_genericstandalone_mon_bussynchronizer63_starter | main_genericstandalone_mon_bussynchronizer63_pong_o) | main_genericstandalone_mon_bussynchronizer63_done);
assign main_genericstandalone_mon_bussynchronizer63_pong_i = main_genericstandalone_mon_bussynchronizer63_ping_o1;
assign main_genericstandalone_mon_bussynchronizer63_ping_o0 = (main_genericstandalone_mon_bussynchronizer63_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer63_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer63_pong_o = (main_genericstandalone_mon_bussynchronizer63_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer63_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer63_done = (main_genericstandalone_mon_bussynchronizer63_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer64_wait = (~main_genericstandalone_mon_bussynchronizer64_ping_i);
assign main_genericstandalone_mon_bussynchronizer64_ping_i = ((main_genericstandalone_mon_bussynchronizer64_starter | main_genericstandalone_mon_bussynchronizer64_pong_o) | main_genericstandalone_mon_bussynchronizer64_done);
assign main_genericstandalone_mon_bussynchronizer64_pong_i = main_genericstandalone_mon_bussynchronizer64_ping_o1;
assign main_genericstandalone_mon_bussynchronizer64_ping_o0 = (main_genericstandalone_mon_bussynchronizer64_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer64_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer64_pong_o = (main_genericstandalone_mon_bussynchronizer64_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer64_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer64_done = (main_genericstandalone_mon_bussynchronizer64_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer65_wait = (~main_genericstandalone_mon_bussynchronizer65_ping_i);
assign main_genericstandalone_mon_bussynchronizer65_ping_i = ((main_genericstandalone_mon_bussynchronizer65_starter | main_genericstandalone_mon_bussynchronizer65_pong_o) | main_genericstandalone_mon_bussynchronizer65_done);
assign main_genericstandalone_mon_bussynchronizer65_pong_i = main_genericstandalone_mon_bussynchronizer65_ping_o1;
assign main_genericstandalone_mon_bussynchronizer65_ping_o0 = (main_genericstandalone_mon_bussynchronizer65_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer65_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer65_pong_o = (main_genericstandalone_mon_bussynchronizer65_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer65_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer65_done = (main_genericstandalone_mon_bussynchronizer65_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer66_wait = (~main_genericstandalone_mon_bussynchronizer66_ping_i);
assign main_genericstandalone_mon_bussynchronizer66_ping_i = ((main_genericstandalone_mon_bussynchronizer66_starter | main_genericstandalone_mon_bussynchronizer66_pong_o) | main_genericstandalone_mon_bussynchronizer66_done);
assign main_genericstandalone_mon_bussynchronizer66_pong_i = main_genericstandalone_mon_bussynchronizer66_ping_o1;
assign main_genericstandalone_mon_bussynchronizer66_ping_o0 = (main_genericstandalone_mon_bussynchronizer66_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer66_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer66_pong_o = (main_genericstandalone_mon_bussynchronizer66_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer66_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer66_done = (main_genericstandalone_mon_bussynchronizer66_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer67_wait = (~main_genericstandalone_mon_bussynchronizer67_ping_i);
assign main_genericstandalone_mon_bussynchronizer67_ping_i = ((main_genericstandalone_mon_bussynchronizer67_starter | main_genericstandalone_mon_bussynchronizer67_pong_o) | main_genericstandalone_mon_bussynchronizer67_done);
assign main_genericstandalone_mon_bussynchronizer67_pong_i = main_genericstandalone_mon_bussynchronizer67_ping_o1;
assign main_genericstandalone_mon_bussynchronizer67_ping_o0 = (main_genericstandalone_mon_bussynchronizer67_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer67_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer67_pong_o = (main_genericstandalone_mon_bussynchronizer67_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer67_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer67_done = (main_genericstandalone_mon_bussynchronizer67_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer68_wait = (~main_genericstandalone_mon_bussynchronizer68_ping_i);
assign main_genericstandalone_mon_bussynchronizer68_ping_i = ((main_genericstandalone_mon_bussynchronizer68_starter | main_genericstandalone_mon_bussynchronizer68_pong_o) | main_genericstandalone_mon_bussynchronizer68_done);
assign main_genericstandalone_mon_bussynchronizer68_pong_i = main_genericstandalone_mon_bussynchronizer68_ping_o1;
assign main_genericstandalone_mon_bussynchronizer68_ping_o0 = (main_genericstandalone_mon_bussynchronizer68_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer68_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer68_pong_o = (main_genericstandalone_mon_bussynchronizer68_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer68_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer68_done = (main_genericstandalone_mon_bussynchronizer68_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer69_wait = (~main_genericstandalone_mon_bussynchronizer69_ping_i);
assign main_genericstandalone_mon_bussynchronizer69_ping_i = ((main_genericstandalone_mon_bussynchronizer69_starter | main_genericstandalone_mon_bussynchronizer69_pong_o) | main_genericstandalone_mon_bussynchronizer69_done);
assign main_genericstandalone_mon_bussynchronizer69_pong_i = main_genericstandalone_mon_bussynchronizer69_ping_o1;
assign main_genericstandalone_mon_bussynchronizer69_ping_o0 = (main_genericstandalone_mon_bussynchronizer69_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer69_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer69_pong_o = (main_genericstandalone_mon_bussynchronizer69_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer69_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer69_done = (main_genericstandalone_mon_bussynchronizer69_count == 1'd0);
assign main_genericstandalone_mon_bussynchronizer70_wait = (~main_genericstandalone_mon_bussynchronizer70_ping_i);
assign main_genericstandalone_mon_bussynchronizer70_ping_i = ((main_genericstandalone_mon_bussynchronizer70_starter | main_genericstandalone_mon_bussynchronizer70_pong_o) | main_genericstandalone_mon_bussynchronizer70_done);
assign main_genericstandalone_mon_bussynchronizer70_pong_i = main_genericstandalone_mon_bussynchronizer70_ping_o1;
assign main_genericstandalone_mon_bussynchronizer70_ping_o0 = (main_genericstandalone_mon_bussynchronizer70_ping_toggle_o ^ main_genericstandalone_mon_bussynchronizer70_ping_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer70_pong_o = (main_genericstandalone_mon_bussynchronizer70_pong_toggle_o ^ main_genericstandalone_mon_bussynchronizer70_pong_toggle_o_r);
assign main_genericstandalone_mon_bussynchronizer70_done = (main_genericstandalone_mon_bussynchronizer70_count == 1'd0);
assign main_genericstandalone_inj_value_w = builder_comb_rhs_self17;
assign main_genericstandalone_rtio_analyzer_fifo_sink_stb = main_genericstandalone_rtio_analyzer_message_encoder_source_stb;
assign main_genericstandalone_rtio_analyzer_message_encoder_source_ack = main_genericstandalone_rtio_analyzer_fifo_sink_ack;
assign main_genericstandalone_rtio_analyzer_fifo_sink_last = main_genericstandalone_rtio_analyzer_message_encoder_source_last;
assign main_genericstandalone_rtio_analyzer_fifo_sink_eop = main_genericstandalone_rtio_analyzer_message_encoder_source_eop;
assign main_genericstandalone_rtio_analyzer_fifo_sink_payload_data = main_genericstandalone_rtio_analyzer_message_encoder_source_payload_data;
assign main_genericstandalone_rtio_analyzer_converter_sink_stb = main_genericstandalone_rtio_analyzer_fifo_source_stb;
assign main_genericstandalone_rtio_analyzer_fifo_source_ack = main_genericstandalone_rtio_analyzer_converter_sink_ack;
assign main_genericstandalone_rtio_analyzer_converter_sink_last = main_genericstandalone_rtio_analyzer_fifo_source_last;
assign main_genericstandalone_rtio_analyzer_converter_sink_eop = main_genericstandalone_rtio_analyzer_fifo_source_eop;
assign main_genericstandalone_rtio_analyzer_converter_sink_payload_data = main_genericstandalone_rtio_analyzer_fifo_source_payload_data;
assign main_genericstandalone_rtio_analyzer_dma_sink_stb = main_genericstandalone_rtio_analyzer_converter_source_stb;
assign main_genericstandalone_rtio_analyzer_converter_source_ack = main_genericstandalone_rtio_analyzer_dma_sink_ack;
assign main_genericstandalone_rtio_analyzer_dma_sink_last = main_genericstandalone_rtio_analyzer_converter_source_last;
assign main_genericstandalone_rtio_analyzer_dma_sink_eop = main_genericstandalone_rtio_analyzer_converter_source_eop;
assign main_genericstandalone_rtio_analyzer_dma_sink_payload_data = main_genericstandalone_rtio_analyzer_converter_source_payload_data;
assign main_genericstandalone_rtio_analyzer_dma_sink_payload_valid_token_count = main_genericstandalone_rtio_analyzer_converter_source_payload_valid_token_count;

// synthesis translate_off
reg dummy_d_212;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_analyzer_message_encoder_read_done <= 1'd0;
	main_genericstandalone_rtio_analyzer_message_encoder_read_overflow <= 1'd0;
	if ((main_genericstandalone_rtio_analyzer_message_encoder_read_wait_event_r & (~main_genericstandalone_rtio_core_cri_i_status[2]))) begin
		if ((~main_genericstandalone_rtio_core_cri_i_status[0])) begin
			main_genericstandalone_rtio_analyzer_message_encoder_read_done <= 1'd1;
		end
		if (main_genericstandalone_rtio_core_cri_i_status[1]) begin
			main_genericstandalone_rtio_analyzer_message_encoder_read_overflow <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_212 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_analyzer_message_encoder_input_output_channel = main_genericstandalone_rtio_core_cri_chan_sel;
assign main_genericstandalone_rtio_analyzer_message_encoder_input_output_address_padding = main_genericstandalone_rtio_core_cri_o_address;
assign main_genericstandalone_rtio_analyzer_message_encoder_input_output_rtio_counter = main_genericstandalone_full_ts;

// synthesis translate_off
reg dummy_d_213;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_analyzer_message_encoder_input_output_message_type <= 2'd0;
	main_genericstandalone_rtio_analyzer_message_encoder_input_output_timestamp <= 64'd0;
	main_genericstandalone_rtio_analyzer_message_encoder_input_output_data <= 64'd0;
	if ((main_genericstandalone_rtio_core_cri_cmd == 1'd1)) begin
		main_genericstandalone_rtio_analyzer_message_encoder_input_output_message_type <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_input_output_timestamp <= main_genericstandalone_rtio_core_cri_o_timestamp;
		main_genericstandalone_rtio_analyzer_message_encoder_input_output_data <= main_genericstandalone_rtio_core_cri_o_data;
	end else begin
		main_genericstandalone_rtio_analyzer_message_encoder_input_output_message_type <= 1'd1;
		main_genericstandalone_rtio_analyzer_message_encoder_input_output_timestamp <= main_genericstandalone_rtio_core_cri_i_timestamp;
		main_genericstandalone_rtio_analyzer_message_encoder_input_output_data <= main_genericstandalone_rtio_core_cri_i_data;
	end
// synthesis translate_off
	dummy_d_213 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_analyzer_message_encoder_input_output_stb = ((main_genericstandalone_rtio_core_cri_cmd == 1'd1) | main_genericstandalone_rtio_analyzer_message_encoder_read_done);
assign main_genericstandalone_rtio_analyzer_message_encoder_exception_message_type = 2'd2;
assign main_genericstandalone_rtio_analyzer_message_encoder_exception_channel = main_genericstandalone_rtio_core_cri_chan_sel;
assign main_genericstandalone_rtio_analyzer_message_encoder_exception_rtio_counter = main_genericstandalone_full_ts;

// synthesis translate_off
reg dummy_d_214;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_analyzer_message_encoder_exception_stb <= 1'd0;
	main_genericstandalone_rtio_analyzer_message_encoder_exception_exception_type <= 8'd0;
	if ((main_genericstandalone_rtio_analyzer_message_encoder_just_written & main_genericstandalone_rtio_core_cri_o_status[1])) begin
		main_genericstandalone_rtio_analyzer_message_encoder_exception_stb <= 1'd1;
		main_genericstandalone_rtio_analyzer_message_encoder_exception_exception_type <= 5'd20;
	end
	if (main_genericstandalone_rtio_analyzer_message_encoder_read_overflow) begin
		main_genericstandalone_rtio_analyzer_message_encoder_exception_stb <= 1'd1;
		main_genericstandalone_rtio_analyzer_message_encoder_exception_exception_type <= 6'd33;
	end
// synthesis translate_off
	dummy_d_214 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_analyzer_message_encoder_stopped_message_type = 2'd3;
assign main_genericstandalone_rtio_analyzer_message_encoder_stopped_rtio_counter = main_genericstandalone_full_ts;
assign main_genericstandalone_rtio_analyzer_fifo_syncfifo_din = {main_genericstandalone_rtio_analyzer_fifo_fifo_in_eop, main_genericstandalone_rtio_analyzer_fifo_fifo_in_payload_data};
assign {main_genericstandalone_rtio_analyzer_fifo_fifo_out_eop, main_genericstandalone_rtio_analyzer_fifo_fifo_out_payload_data} = main_genericstandalone_rtio_analyzer_fifo_syncfifo_dout;
assign main_genericstandalone_rtio_analyzer_fifo_sink_ack = main_genericstandalone_rtio_analyzer_fifo_syncfifo_writable;
assign main_genericstandalone_rtio_analyzer_fifo_syncfifo_we = main_genericstandalone_rtio_analyzer_fifo_sink_stb;
assign main_genericstandalone_rtio_analyzer_fifo_fifo_in_eop = main_genericstandalone_rtio_analyzer_fifo_sink_eop;
assign main_genericstandalone_rtio_analyzer_fifo_fifo_in_payload_data = main_genericstandalone_rtio_analyzer_fifo_sink_payload_data;
assign main_genericstandalone_rtio_analyzer_fifo_source_eop = main_genericstandalone_rtio_analyzer_fifo_fifo_out_eop;
assign main_genericstandalone_rtio_analyzer_fifo_source_payload_data = main_genericstandalone_rtio_analyzer_fifo_fifo_out_payload_data;

// synthesis translate_off
reg dummy_d_215;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_analyzer_fifo_re <= 1'd0;
	main_genericstandalone_rtio_analyzer_fifo_re <= main_genericstandalone_rtio_analyzer_fifo_source_ack;
	main_genericstandalone_rtio_analyzer_fifo_re <= (main_genericstandalone_rtio_analyzer_fifo_source_stb & main_genericstandalone_rtio_analyzer_fifo_source_ack);
// synthesis translate_off
	dummy_d_215 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_analyzer_fifo_do_write = (main_genericstandalone_rtio_analyzer_fifo_syncfifo_we & main_genericstandalone_rtio_analyzer_fifo_syncfifo_writable);
assign main_genericstandalone_rtio_analyzer_fifo_do_read1 = (main_genericstandalone_rtio_analyzer_fifo_re & main_genericstandalone_rtio_analyzer_fifo_readable);
assign main_genericstandalone_rtio_analyzer_fifo_has_pending_eop = (main_genericstandalone_rtio_analyzer_fifo_eop_count_next != 1'd0);

// synthesis translate_off
reg dummy_d_216;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_analyzer_fifo_eop_count_next <= 8'd0;
	main_genericstandalone_rtio_analyzer_fifo_eop_count_next <= main_genericstandalone_rtio_analyzer_fifo_eop_count;
	if ((main_genericstandalone_rtio_analyzer_fifo_fifo_in_eop & main_genericstandalone_rtio_analyzer_fifo_do_write)) begin
		if ((~(main_genericstandalone_rtio_analyzer_fifo_fifo_out_eop & main_genericstandalone_rtio_analyzer_fifo_do_read1))) begin
			main_genericstandalone_rtio_analyzer_fifo_eop_count_next <= (main_genericstandalone_rtio_analyzer_fifo_eop_count + 1'd1);
		end
	end else begin
		if ((main_genericstandalone_rtio_analyzer_fifo_fifo_out_eop & main_genericstandalone_rtio_analyzer_fifo_do_read1)) begin
			main_genericstandalone_rtio_analyzer_fifo_eop_count_next <= (main_genericstandalone_rtio_analyzer_fifo_eop_count - 1'd1);
		end
	end
// synthesis translate_off
	dummy_d_216 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_analyzer_fifo_source_last = ((main_genericstandalone_rtio_analyzer_fifo_transfer_count == 1'd0) | main_genericstandalone_rtio_analyzer_fifo_fifo_out_eop);

// synthesis translate_off
reg dummy_d_217;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_analyzer_fifo_source_stb <= 1'd0;
	main_genericstandalone_rtio_analyzer_fifo_source_stb <= main_genericstandalone_rtio_analyzer_fifo_readable;
	main_genericstandalone_rtio_analyzer_fifo_source_stb <= (main_genericstandalone_rtio_analyzer_fifo_readable & (main_genericstandalone_rtio_analyzer_fifo_almost_full | main_genericstandalone_rtio_analyzer_fifo_activated));
// synthesis translate_off
	dummy_d_217 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_analyzer_fifo_transfer_count_ce = main_genericstandalone_rtio_analyzer_fifo_do_read1;
assign main_genericstandalone_rtio_analyzer_fifo_transfer_count_rst = (main_genericstandalone_rtio_analyzer_fifo_do_read1 & main_genericstandalone_rtio_analyzer_fifo_source_last);
assign main_genericstandalone_rtio_analyzer_fifo_syncfifo_re = (main_genericstandalone_rtio_analyzer_fifo_syncfifo_readable & ((~main_genericstandalone_rtio_analyzer_fifo_readable) | main_genericstandalone_rtio_analyzer_fifo_re));
assign main_genericstandalone_rtio_analyzer_fifo_level1 = (main_genericstandalone_rtio_analyzer_fifo_level0 + main_genericstandalone_rtio_analyzer_fifo_readable);
assign main_genericstandalone_rtio_analyzer_fifo_almost_full = (main_genericstandalone_rtio_analyzer_fifo_level1 >= 7'd64);

// synthesis translate_off
reg dummy_d_218;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_analyzer_fifo_wrport_adr <= 7'd0;
	if (main_genericstandalone_rtio_analyzer_fifo_replace) begin
		main_genericstandalone_rtio_analyzer_fifo_wrport_adr <= (main_genericstandalone_rtio_analyzer_fifo_produce - 1'd1);
	end else begin
		main_genericstandalone_rtio_analyzer_fifo_wrport_adr <= main_genericstandalone_rtio_analyzer_fifo_produce;
	end
// synthesis translate_off
	dummy_d_218 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_analyzer_fifo_wrport_dat_w = main_genericstandalone_rtio_analyzer_fifo_syncfifo_din;
assign main_genericstandalone_rtio_analyzer_fifo_wrport_we = (main_genericstandalone_rtio_analyzer_fifo_syncfifo_we & (main_genericstandalone_rtio_analyzer_fifo_syncfifo_writable | main_genericstandalone_rtio_analyzer_fifo_replace));
assign main_genericstandalone_rtio_analyzer_fifo_do_read0 = (main_genericstandalone_rtio_analyzer_fifo_syncfifo_readable & main_genericstandalone_rtio_analyzer_fifo_syncfifo_re);
assign main_genericstandalone_rtio_analyzer_fifo_rdport_adr = main_genericstandalone_rtio_analyzer_fifo_consume;
assign main_genericstandalone_rtio_analyzer_fifo_syncfifo_dout = main_genericstandalone_rtio_analyzer_fifo_rdport_dat_r;
assign main_genericstandalone_rtio_analyzer_fifo_rdport_re = main_genericstandalone_rtio_analyzer_fifo_do_read0;
assign main_genericstandalone_rtio_analyzer_fifo_syncfifo_writable = (main_genericstandalone_rtio_analyzer_fifo_level0 != 8'd128);
assign main_genericstandalone_rtio_analyzer_fifo_syncfifo_readable = (main_genericstandalone_rtio_analyzer_fifo_level0 != 1'd0);
assign main_genericstandalone_rtio_analyzer_converter_last = (main_genericstandalone_rtio_analyzer_converter_mux == 1'd1);
assign main_genericstandalone_rtio_analyzer_converter_source_stb = main_genericstandalone_rtio_analyzer_converter_sink_stb;
assign main_genericstandalone_rtio_analyzer_converter_source_eop = (main_genericstandalone_rtio_analyzer_converter_sink_eop & main_genericstandalone_rtio_analyzer_converter_last);
assign main_genericstandalone_rtio_analyzer_converter_source_last = (main_genericstandalone_rtio_analyzer_converter_sink_last & main_genericstandalone_rtio_analyzer_converter_last);
assign main_genericstandalone_rtio_analyzer_converter_sink_ack = (main_genericstandalone_rtio_analyzer_converter_last & main_genericstandalone_rtio_analyzer_converter_source_ack);

// synthesis translate_off
reg dummy_d_219;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rtio_analyzer_converter_source_payload_data <= 128'd0;
	case (main_genericstandalone_rtio_analyzer_converter_mux)
		1'd0: begin
			main_genericstandalone_rtio_analyzer_converter_source_payload_data <= main_genericstandalone_rtio_analyzer_converter_sink_payload_data[255:128];
		end
		default: begin
			main_genericstandalone_rtio_analyzer_converter_source_payload_data <= main_genericstandalone_rtio_analyzer_converter_sink_payload_data[127:0];
		end
	endcase
// synthesis translate_off
	dummy_d_219 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rtio_analyzer_converter_source_payload_valid_token_count = main_genericstandalone_rtio_analyzer_converter_last;
assign main_genericstandalone_interface1_bus_cyc = main_genericstandalone_rtio_analyzer_dma_sink_stb;
assign main_genericstandalone_interface1_bus_stb = main_genericstandalone_rtio_analyzer_dma_sink_stb;
assign main_genericstandalone_interface1_bus_cti = (main_genericstandalone_rtio_analyzer_dma_sink_last ? 3'd7 : 2'd2);
assign main_genericstandalone_rtio_analyzer_dma_sink_ack = main_genericstandalone_interface1_bus_ack;
assign main_genericstandalone_interface1_bus_we = 1'd1;
assign main_genericstandalone_interface1_bus_dat_w = {{builder_slice_proxy31[7:0], builder_slice_proxy30[15:8], builder_slice_proxy29[23:16], builder_slice_proxy28[31:24], builder_slice_proxy27[39:32], builder_slice_proxy26[47:40], builder_slice_proxy25[55:48], builder_slice_proxy24[63:56]}, {builder_slice_proxy23[7:0], builder_slice_proxy22[15:8], builder_slice_proxy21[23:16], builder_slice_proxy20[31:24], builder_slice_proxy19[39:32], builder_slice_proxy18[47:40], builder_slice_proxy17[55:48], builder_slice_proxy16[63:56]}};
assign main_genericstandalone_interface1_bus_sel = 16'd65535;
assign main_genericstandalone_rtio_analyzer_dma_status = (main_genericstandalone_rtio_analyzer_dma_message_count <<< 3'd5);
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr = builder_comb_rhs_self56;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_w = builder_comb_rhs_self57;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel = builder_comb_rhs_self58;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cyc = builder_comb_rhs_self59;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_stb = builder_comb_rhs_self60;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_we = builder_comb_rhs_self61;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cti = builder_comb_rhs_self62;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_bte = builder_comb_rhs_self63;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_r = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r;
assign main_genericstandalone_kernel_cpu_wb_sdram_dat_r = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_ack = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack & (builder_sdram_cpulevel_arbiter_grant == 1'd0));
assign main_genericstandalone_kernel_cpu_wb_sdram_ack = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack & (builder_sdram_cpulevel_arbiter_grant == 1'd1));
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_err = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_err & (builder_sdram_cpulevel_arbiter_grant == 1'd0));
assign main_genericstandalone_kernel_cpu_wb_sdram_err = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_err & (builder_sdram_cpulevel_arbiter_grant == 1'd1));
assign builder_sdram_cpulevel_arbiter_request = {(main_genericstandalone_kernel_cpu_wb_sdram_cyc & (~(main_genericstandalone_kernel_cpu_wb_sdram_ack & (main_genericstandalone_kernel_cpu_wb_sdram_cti != 2'd2)))), (main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cyc & (~(main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_ack & (main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cti != 2'd2))))};
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr = builder_comb_rhs_self64;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_w = builder_comb_rhs_self65;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_sel = builder_comb_rhs_self66;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cyc = builder_comb_rhs_self67;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_stb = builder_comb_rhs_self68;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_we = builder_comb_rhs_self69;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti = builder_comb_rhs_self70;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_bte = builder_comb_rhs_self71;
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r;
assign main_genericstandalone_interface0_bus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r;
assign main_genericstandalone_interface1_bus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 1'd0));
assign main_genericstandalone_interface0_bus_ack = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 1'd1));
assign main_genericstandalone_interface1_bus_ack = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 2'd2));
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_err = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 1'd0));
assign main_genericstandalone_interface0_bus_err = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 1'd1));
assign main_genericstandalone_interface1_bus_err = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 2'd2));
assign builder_sdram_native_arbiter_request = {(main_genericstandalone_interface1_bus_cyc & (~(main_genericstandalone_interface1_bus_ack & (main_genericstandalone_interface1_bus_cti != 2'd2)))), (main_genericstandalone_interface0_bus_cyc & (~(main_genericstandalone_interface0_bus_ack & (main_genericstandalone_interface0_bus_cti != 2'd2)))), (main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc & (~(main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack & (main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cti != 2'd2))))};
assign builder_genericstandalone_shared_adr = builder_comb_rhs_self72;
assign builder_genericstandalone_shared_dat_w = builder_comb_rhs_self73;
assign builder_genericstandalone_shared_sel = builder_comb_rhs_self74;
assign builder_genericstandalone_shared_cyc = builder_comb_rhs_self75;
assign builder_genericstandalone_shared_stb = builder_comb_rhs_self76;
assign builder_genericstandalone_shared_we = builder_comb_rhs_self77;
assign builder_genericstandalone_shared_cti = builder_comb_rhs_self78;
assign builder_genericstandalone_shared_bte = builder_comb_rhs_self79;
assign main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_r = builder_genericstandalone_shared_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_r = builder_genericstandalone_shared_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_ibus_ack = (builder_genericstandalone_shared_ack & (builder_genericstandalone_grant == 1'd0));
assign main_genericstandalone_genericstandalone_genericstandalone_dbus_ack = (builder_genericstandalone_shared_ack & (builder_genericstandalone_grant == 1'd1));
assign main_genericstandalone_genericstandalone_genericstandalone_ibus_err = (builder_genericstandalone_shared_err & (builder_genericstandalone_grant == 1'd0));
assign main_genericstandalone_genericstandalone_genericstandalone_dbus_err = (builder_genericstandalone_shared_err & (builder_genericstandalone_grant == 1'd1));
assign builder_genericstandalone_request = {(main_genericstandalone_genericstandalone_genericstandalone_dbus_cyc & (~(main_genericstandalone_genericstandalone_genericstandalone_dbus_ack & (main_genericstandalone_genericstandalone_genericstandalone_dbus_cti != 2'd2)))), (main_genericstandalone_genericstandalone_genericstandalone_ibus_cyc & (~(main_genericstandalone_genericstandalone_genericstandalone_ibus_ack & (main_genericstandalone_genericstandalone_genericstandalone_ibus_cti != 2'd2))))};

// synthesis translate_off
reg dummy_d_220;
// synthesis translate_on
always @(*) begin
	builder_genericstandalone_slave_sel <= 6'd0;
	builder_genericstandalone_slave_sel[0] <= (((1'd1 & (~builder_genericstandalone_shared_adr[26])) & (~builder_genericstandalone_shared_adr[27])) & builder_genericstandalone_shared_adr[25]);
	builder_genericstandalone_slave_sel[1] <= (((1'd1 & (~builder_genericstandalone_shared_adr[25])) & builder_genericstandalone_shared_adr[26]) & builder_genericstandalone_shared_adr[27]);
	builder_genericstandalone_slave_sel[2] <= ((1'd1 & (~builder_genericstandalone_shared_adr[26])) & builder_genericstandalone_shared_adr[27]);
	builder_genericstandalone_slave_sel[3] <= (((1'd1 & (~builder_genericstandalone_shared_adr[25])) & (~builder_genericstandalone_shared_adr[26])) & (~builder_genericstandalone_shared_adr[27]));
	builder_genericstandalone_slave_sel[4] <= ((1'd1 & (~builder_genericstandalone_shared_adr[27])) & builder_genericstandalone_shared_adr[26]);
	builder_genericstandalone_slave_sel[5] <= (((1'd1 & builder_genericstandalone_shared_adr[25]) & builder_genericstandalone_shared_adr[26]) & builder_genericstandalone_shared_adr[27]);
// synthesis translate_off
	dummy_d_220 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_genericstandalone_spiflash_bus_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_genericstandalone_spiflash_bus_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_genericstandalone_spiflash_bus_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_genericstandalone_spiflash_bus_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_genericstandalone_spiflash_bus_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_genericstandalone_spiflash_bus_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_genericstandalone_spiflash_bus_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_bus_bus_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_bus_bus_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_bus_bus_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_bus_bus_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_bus_bus_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_bus_bus_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_bus_bus_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_mailbox_i1_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_mailbox_i1_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_mailbox_i1_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_mailbox_i1_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_mailbox_i1_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_mailbox_i1_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_mailbox_i1_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[0]);
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[1]);
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[2]);
assign main_genericstandalone_genericstandalone_spiflash_bus_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[3]);
assign main_genericstandalone_bus_bus_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[4]);
assign main_genericstandalone_mailbox_i1_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[5]);
assign builder_genericstandalone_shared_ack = (((((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack | main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack) | main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_ack) | main_genericstandalone_genericstandalone_spiflash_bus_ack) | main_genericstandalone_bus_bus_ack) | main_genericstandalone_mailbox_i1_ack);
assign builder_genericstandalone_shared_err = (((((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_err | main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_err) | main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_err) | main_genericstandalone_genericstandalone_spiflash_bus_err) | main_genericstandalone_bus_bus_err) | main_genericstandalone_mailbox_i1_err);
assign builder_genericstandalone_shared_dat_r = (((((({64{builder_genericstandalone_slave_sel_r[0]}} & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_r) | ({64{builder_genericstandalone_slave_sel_r[1]}} & main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_r)) | ({64{builder_genericstandalone_slave_sel_r[2]}} & main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_r)) | ({64{builder_genericstandalone_slave_sel_r[3]}} & main_genericstandalone_genericstandalone_spiflash_bus_dat_r)) | ({64{builder_genericstandalone_slave_sel_r[4]}} & main_genericstandalone_bus_bus_dat_r)) | ({64{builder_genericstandalone_slave_sel_r[5]}} & main_genericstandalone_mailbox_i1_dat_r));
assign builder_genericstandalone_csrbank0_sel = (builder_genericstandalone_interface0_bank_bus_adr[13:8] == 3'd6);
assign builder_genericstandalone_csrbank0_switch_done_r = builder_genericstandalone_interface0_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank0_switch_done_re = ((builder_genericstandalone_csrbank0_sel & builder_genericstandalone_interface0_bank_bus_we) & (builder_genericstandalone_interface0_bank_bus_adr[0] == 1'd0));
assign builder_genericstandalone_csrbank0_clock_sel0_r = builder_genericstandalone_interface0_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank0_clock_sel0_re = ((builder_genericstandalone_csrbank0_sel & builder_genericstandalone_interface0_bank_bus_we) & (builder_genericstandalone_interface0_bank_bus_adr[0] == 1'd1));
assign builder_genericstandalone_csrbank0_switch_done_w = main_genericstandalone_genericstandalone_crg_status;
assign main_genericstandalone_rtiosyscrg_storage = main_genericstandalone_rtiosyscrg_storage_full;
assign builder_genericstandalone_csrbank0_clock_sel0_w = main_genericstandalone_rtiosyscrg_storage_full;
assign builder_genericstandalone_csrbank1_sel = (builder_genericstandalone_interface1_bank_bus_adr[13:8] == 3'd7);
assign builder_genericstandalone_csrbank1_dly_sel0_r = builder_genericstandalone_interface1_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank1_dly_sel0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[1:0] == 1'd0));
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_r = builder_genericstandalone_interface1_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[1:0] == 1'd1));
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_r = builder_genericstandalone_interface1_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[1:0] == 2'd2));
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_r = builder_genericstandalone_interface1_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[1:0] == 2'd3));
assign main_genericstandalone_genericstandalone_ddrphy_storage = main_genericstandalone_genericstandalone_ddrphy_storage_full[1:0];
assign builder_genericstandalone_csrbank1_dly_sel0_w = main_genericstandalone_genericstandalone_ddrphy_storage_full[1:0];
assign builder_genericstandalone_csrbank2_sel = (builder_genericstandalone_interface2_bank_bus_adr[13:8] == 3'd4);
assign builder_genericstandalone_csrbank2_control0_r = builder_genericstandalone_interface2_bank_bus_dat_w[3:0];
assign builder_genericstandalone_csrbank2_control0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 1'd0));
assign builder_genericstandalone_csrbank2_pi0_command0_r = builder_genericstandalone_interface2_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank2_pi0_command0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 1'd1));
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 2'd2));
assign builder_genericstandalone_csrbank2_pi0_address1_r = builder_genericstandalone_interface2_bank_bus_dat_w[6:0];
assign builder_genericstandalone_csrbank2_pi0_address1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 2'd3));
assign builder_genericstandalone_csrbank2_pi0_address0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_address0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 3'd4));
assign builder_genericstandalone_csrbank2_pi0_baddress0_r = builder_genericstandalone_interface2_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank2_pi0_baddress0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 3'd5));
assign builder_genericstandalone_csrbank2_pi0_wrdata3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_wrdata3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 3'd6));
assign builder_genericstandalone_csrbank2_pi0_wrdata2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_wrdata2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 3'd7));
assign builder_genericstandalone_csrbank2_pi0_wrdata1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_wrdata1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 4'd8));
assign builder_genericstandalone_csrbank2_pi0_wrdata0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_wrdata0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 4'd9));
assign builder_genericstandalone_csrbank2_pi0_rddata3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_rddata3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 4'd10));
assign builder_genericstandalone_csrbank2_pi0_rddata2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_rddata2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 4'd11));
assign builder_genericstandalone_csrbank2_pi0_rddata1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_rddata1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 4'd12));
assign builder_genericstandalone_csrbank2_pi0_rddata0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi0_rddata0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 4'd13));
assign builder_genericstandalone_csrbank2_pi1_command0_r = builder_genericstandalone_interface2_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank2_pi1_command0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 4'd14));
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 4'd15));
assign builder_genericstandalone_csrbank2_pi1_address1_r = builder_genericstandalone_interface2_bank_bus_dat_w[6:0];
assign builder_genericstandalone_csrbank2_pi1_address1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd16));
assign builder_genericstandalone_csrbank2_pi1_address0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_address0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd17));
assign builder_genericstandalone_csrbank2_pi1_baddress0_r = builder_genericstandalone_interface2_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank2_pi1_baddress0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd18));
assign builder_genericstandalone_csrbank2_pi1_wrdata3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_wrdata3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd19));
assign builder_genericstandalone_csrbank2_pi1_wrdata2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_wrdata2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd20));
assign builder_genericstandalone_csrbank2_pi1_wrdata1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_wrdata1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd21));
assign builder_genericstandalone_csrbank2_pi1_wrdata0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_wrdata0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd22));
assign builder_genericstandalone_csrbank2_pi1_rddata3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_rddata3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd23));
assign builder_genericstandalone_csrbank2_pi1_rddata2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_rddata2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd24));
assign builder_genericstandalone_csrbank2_pi1_rddata1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_rddata1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd25));
assign builder_genericstandalone_csrbank2_pi1_rddata0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi1_rddata0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd26));
assign builder_genericstandalone_csrbank2_pi2_command0_r = builder_genericstandalone_interface2_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank2_pi2_command0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd27));
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd28));
assign builder_genericstandalone_csrbank2_pi2_address1_r = builder_genericstandalone_interface2_bank_bus_dat_w[6:0];
assign builder_genericstandalone_csrbank2_pi2_address1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd29));
assign builder_genericstandalone_csrbank2_pi2_address0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_address0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd30));
assign builder_genericstandalone_csrbank2_pi2_baddress0_r = builder_genericstandalone_interface2_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank2_pi2_baddress0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 5'd31));
assign builder_genericstandalone_csrbank2_pi2_wrdata3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_wrdata3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd32));
assign builder_genericstandalone_csrbank2_pi2_wrdata2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_wrdata2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd33));
assign builder_genericstandalone_csrbank2_pi2_wrdata1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_wrdata1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd34));
assign builder_genericstandalone_csrbank2_pi2_wrdata0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_wrdata0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd35));
assign builder_genericstandalone_csrbank2_pi2_rddata3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_rddata3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd36));
assign builder_genericstandalone_csrbank2_pi2_rddata2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_rddata2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd37));
assign builder_genericstandalone_csrbank2_pi2_rddata1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_rddata1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd38));
assign builder_genericstandalone_csrbank2_pi2_rddata0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi2_rddata0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd39));
assign builder_genericstandalone_csrbank2_pi3_command0_r = builder_genericstandalone_interface2_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank2_pi3_command0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd40));
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd41));
assign builder_genericstandalone_csrbank2_pi3_address1_r = builder_genericstandalone_interface2_bank_bus_dat_w[6:0];
assign builder_genericstandalone_csrbank2_pi3_address1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd42));
assign builder_genericstandalone_csrbank2_pi3_address0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_address0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd43));
assign builder_genericstandalone_csrbank2_pi3_baddress0_r = builder_genericstandalone_interface2_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank2_pi3_baddress0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd44));
assign builder_genericstandalone_csrbank2_pi3_wrdata3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_wrdata3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd45));
assign builder_genericstandalone_csrbank2_pi3_wrdata2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_wrdata2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd46));
assign builder_genericstandalone_csrbank2_pi3_wrdata1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_wrdata1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd47));
assign builder_genericstandalone_csrbank2_pi3_wrdata0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_wrdata0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd48));
assign builder_genericstandalone_csrbank2_pi3_rddata3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_rddata3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd49));
assign builder_genericstandalone_csrbank2_pi3_rddata2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_rddata2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd50));
assign builder_genericstandalone_csrbank2_pi3_rddata1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_rddata1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd51));
assign builder_genericstandalone_csrbank2_pi3_rddata0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_pi3_rddata0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[5:0] == 6'd52));
assign main_genericstandalone_genericstandalone_genericstandalone_storage = main_genericstandalone_genericstandalone_genericstandalone_storage_full[3:0];
assign builder_genericstandalone_csrbank2_control0_w = main_genericstandalone_genericstandalone_genericstandalone_storage_full[3:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full[5:0];
assign builder_genericstandalone_csrbank2_pi0_command0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full[5:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[14:0];
assign builder_genericstandalone_csrbank2_pi0_address1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[14:8];
assign builder_genericstandalone_csrbank2_pi0_address0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full[2:0];
assign builder_genericstandalone_csrbank2_pi0_baddress0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full[2:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[31:0];
assign builder_genericstandalone_csrbank2_pi0_wrdata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[31:24];
assign builder_genericstandalone_csrbank2_pi0_wrdata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[23:16];
assign builder_genericstandalone_csrbank2_pi0_wrdata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[15:8];
assign builder_genericstandalone_csrbank2_pi0_wrdata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[7:0];
assign builder_genericstandalone_csrbank2_pi0_rddata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status[31:24];
assign builder_genericstandalone_csrbank2_pi0_rddata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status[23:16];
assign builder_genericstandalone_csrbank2_pi0_rddata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status[15:8];
assign builder_genericstandalone_csrbank2_pi0_rddata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full[5:0];
assign builder_genericstandalone_csrbank2_pi1_command0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full[5:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[14:0];
assign builder_genericstandalone_csrbank2_pi1_address1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[14:8];
assign builder_genericstandalone_csrbank2_pi1_address0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full[2:0];
assign builder_genericstandalone_csrbank2_pi1_baddress0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full[2:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[31:0];
assign builder_genericstandalone_csrbank2_pi1_wrdata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[31:24];
assign builder_genericstandalone_csrbank2_pi1_wrdata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[23:16];
assign builder_genericstandalone_csrbank2_pi1_wrdata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[15:8];
assign builder_genericstandalone_csrbank2_pi1_wrdata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[7:0];
assign builder_genericstandalone_csrbank2_pi1_rddata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status[31:24];
assign builder_genericstandalone_csrbank2_pi1_rddata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status[23:16];
assign builder_genericstandalone_csrbank2_pi1_rddata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status[15:8];
assign builder_genericstandalone_csrbank2_pi1_rddata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full[5:0];
assign builder_genericstandalone_csrbank2_pi2_command0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full[5:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[14:0];
assign builder_genericstandalone_csrbank2_pi2_address1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[14:8];
assign builder_genericstandalone_csrbank2_pi2_address0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full[2:0];
assign builder_genericstandalone_csrbank2_pi2_baddress0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full[2:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[31:0];
assign builder_genericstandalone_csrbank2_pi2_wrdata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[31:24];
assign builder_genericstandalone_csrbank2_pi2_wrdata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[23:16];
assign builder_genericstandalone_csrbank2_pi2_wrdata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[15:8];
assign builder_genericstandalone_csrbank2_pi2_wrdata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[7:0];
assign builder_genericstandalone_csrbank2_pi2_rddata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status[31:24];
assign builder_genericstandalone_csrbank2_pi2_rddata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status[23:16];
assign builder_genericstandalone_csrbank2_pi2_rddata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status[15:8];
assign builder_genericstandalone_csrbank2_pi2_rddata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full[5:0];
assign builder_genericstandalone_csrbank2_pi3_command0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full[5:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[14:0];
assign builder_genericstandalone_csrbank2_pi3_address1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[14:8];
assign builder_genericstandalone_csrbank2_pi3_address0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full[2:0];
assign builder_genericstandalone_csrbank2_pi3_baddress0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full[2:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[31:0];
assign builder_genericstandalone_csrbank2_pi3_wrdata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[31:24];
assign builder_genericstandalone_csrbank2_pi3_wrdata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[23:16];
assign builder_genericstandalone_csrbank2_pi3_wrdata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[15:8];
assign builder_genericstandalone_csrbank2_pi3_wrdata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[7:0];
assign builder_genericstandalone_csrbank2_pi3_rddata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status[31:24];
assign builder_genericstandalone_csrbank2_pi3_rddata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status[23:16];
assign builder_genericstandalone_csrbank2_pi3_rddata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status[15:8];
assign builder_genericstandalone_csrbank2_pi3_rddata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status[7:0];
assign builder_genericstandalone_csrbank3_sel = (builder_genericstandalone_interface3_bank_bus_adr[13:8] == 4'd14);
assign builder_genericstandalone_csrbank3_out0_r = builder_genericstandalone_interface3_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank3_out0_re = ((builder_genericstandalone_csrbank3_sel & builder_genericstandalone_interface3_bank_bus_we) & (builder_genericstandalone_interface3_bank_bus_adr[0] == 1'd0));
assign main_genericstandalone_error_led_storage = main_genericstandalone_error_led_storage_full;
assign builder_genericstandalone_csrbank3_out0_w = main_genericstandalone_error_led_storage_full;
assign builder_genericstandalone_csrbank4_sel = (builder_genericstandalone_interface4_bank_bus_adr[13:8] == 4'd12);
assign builder_genericstandalone_csrbank4_sram_writer_slot_r = builder_genericstandalone_interface4_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank4_sram_writer_slot_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 1'd0));
assign builder_genericstandalone_csrbank4_sram_writer_length1_r = builder_genericstandalone_interface4_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank4_sram_writer_length1_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 1'd1));
assign builder_genericstandalone_csrbank4_sram_writer_length0_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_sram_writer_length0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 2'd2));
assign builder_genericstandalone_csrbank4_sram_writer_errors3_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_sram_writer_errors3_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 2'd3));
assign builder_genericstandalone_csrbank4_sram_writer_errors2_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_sram_writer_errors2_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 3'd4));
assign builder_genericstandalone_csrbank4_sram_writer_errors1_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_sram_writer_errors1_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 3'd5));
assign builder_genericstandalone_csrbank4_sram_writer_errors0_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_sram_writer_errors0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 3'd6));
assign main_genericstandalone_sram24_status_r = builder_genericstandalone_interface4_bank_bus_dat_w[0];
assign main_genericstandalone_sram23_status_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 3'd7));
assign main_genericstandalone_sram27_pending_r = builder_genericstandalone_interface4_bank_bus_dat_w[0];
assign main_genericstandalone_sram26_pending_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 4'd8));
assign builder_genericstandalone_csrbank4_sram_writer_ev_enable0_r = builder_genericstandalone_interface4_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank4_sram_writer_ev_enable0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 4'd9));
assign main_genericstandalone_start_r = builder_genericstandalone_interface4_bank_bus_dat_w[0];
assign main_genericstandalone_start_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 4'd10));
assign builder_genericstandalone_csrbank4_sram_reader_ready_r = builder_genericstandalone_interface4_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank4_sram_reader_ready_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 4'd11));
assign builder_genericstandalone_csrbank4_sram_reader_slot0_r = builder_genericstandalone_interface4_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank4_sram_reader_slot0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 4'd12));
assign builder_genericstandalone_csrbank4_sram_reader_length1_r = builder_genericstandalone_interface4_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank4_sram_reader_length1_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 4'd13));
assign builder_genericstandalone_csrbank4_sram_reader_length0_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_sram_reader_length0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 4'd14));
assign main_genericstandalone_sram111_status_r = builder_genericstandalone_interface4_bank_bus_dat_w[0];
assign main_genericstandalone_sram110_status_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 4'd15));
assign main_genericstandalone_sram114_pending_r = builder_genericstandalone_interface4_bank_bus_dat_w[0];
assign main_genericstandalone_sram113_pending_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd16));
assign builder_genericstandalone_csrbank4_sram_reader_ev_enable0_r = builder_genericstandalone_interface4_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank4_sram_reader_ev_enable0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd17));
assign builder_genericstandalone_csrbank4_preamble_errors3_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_preamble_errors3_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd18));
assign builder_genericstandalone_csrbank4_preamble_errors2_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_preamble_errors2_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd19));
assign builder_genericstandalone_csrbank4_preamble_errors1_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_preamble_errors1_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd20));
assign builder_genericstandalone_csrbank4_preamble_errors0_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_preamble_errors0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd21));
assign builder_genericstandalone_csrbank4_crc_errors3_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_crc_errors3_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd22));
assign builder_genericstandalone_csrbank4_crc_errors2_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_crc_errors2_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd23));
assign builder_genericstandalone_csrbank4_crc_errors1_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_crc_errors1_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd24));
assign builder_genericstandalone_csrbank4_crc_errors0_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_crc_errors0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[4:0] == 5'd25));
assign builder_genericstandalone_csrbank4_sram_writer_slot_w = main_genericstandalone_sram15_status[1:0];
assign builder_genericstandalone_csrbank4_sram_writer_length1_w = main_genericstandalone_sram16_status[10:8];
assign builder_genericstandalone_csrbank4_sram_writer_length0_w = main_genericstandalone_sram16_status[7:0];
assign builder_genericstandalone_csrbank4_sram_writer_errors3_w = main_genericstandalone_sram17_status[31:24];
assign builder_genericstandalone_csrbank4_sram_writer_errors2_w = main_genericstandalone_sram17_status[23:16];
assign builder_genericstandalone_csrbank4_sram_writer_errors1_w = main_genericstandalone_sram17_status[15:8];
assign builder_genericstandalone_csrbank4_sram_writer_errors0_w = main_genericstandalone_sram17_status[7:0];
assign main_genericstandalone_sram30_storage = main_genericstandalone_sram29_storage_full;
assign builder_genericstandalone_csrbank4_sram_writer_ev_enable0_w = main_genericstandalone_sram29_storage_full;
assign builder_genericstandalone_csrbank4_sram_reader_ready_w = main_genericstandalone_sram98_status;
assign main_genericstandalone_sram100_storage = main_genericstandalone_sram99_storage_full[1:0];
assign builder_genericstandalone_csrbank4_sram_reader_slot0_w = main_genericstandalone_sram99_storage_full[1:0];
assign main_genericstandalone_sram103_storage = main_genericstandalone_sram102_storage_full[10:0];
assign builder_genericstandalone_csrbank4_sram_reader_length1_w = main_genericstandalone_sram102_storage_full[10:8];
assign builder_genericstandalone_csrbank4_sram_reader_length0_w = main_genericstandalone_sram102_storage_full[7:0];
assign main_genericstandalone_sram117_storage = main_genericstandalone_sram116_storage_full;
assign builder_genericstandalone_csrbank4_sram_reader_ev_enable0_w = main_genericstandalone_sram116_storage_full;
assign builder_genericstandalone_csrbank4_preamble_errors3_w = main_genericstandalone_preamble_errors_status[31:24];
assign builder_genericstandalone_csrbank4_preamble_errors2_w = main_genericstandalone_preamble_errors_status[23:16];
assign builder_genericstandalone_csrbank4_preamble_errors1_w = main_genericstandalone_preamble_errors_status[15:8];
assign builder_genericstandalone_csrbank4_preamble_errors0_w = main_genericstandalone_preamble_errors_status[7:0];
assign builder_genericstandalone_csrbank4_crc_errors3_w = main_genericstandalone_crc_errors_status[31:24];
assign builder_genericstandalone_csrbank4_crc_errors2_w = main_genericstandalone_crc_errors_status[23:16];
assign builder_genericstandalone_csrbank4_crc_errors1_w = main_genericstandalone_crc_errors_status[15:8];
assign builder_genericstandalone_csrbank4_crc_errors0_w = main_genericstandalone_crc_errors_status[7:0];
assign builder_genericstandalone_csrbank5_sel = (builder_genericstandalone_interface5_bank_bus_adr[13:8] == 4'd15);
assign builder_genericstandalone_csrbank5_in_r = builder_genericstandalone_interface5_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank5_in_re = ((builder_genericstandalone_csrbank5_sel & builder_genericstandalone_interface5_bank_bus_we) & (builder_genericstandalone_interface5_bank_bus_adr[1:0] == 1'd0));
assign builder_genericstandalone_csrbank5_out0_r = builder_genericstandalone_interface5_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank5_out0_re = ((builder_genericstandalone_csrbank5_sel & builder_genericstandalone_interface5_bank_bus_we) & (builder_genericstandalone_interface5_bank_bus_adr[1:0] == 1'd1));
assign builder_genericstandalone_csrbank5_oe0_r = builder_genericstandalone_interface5_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank5_oe0_re = ((builder_genericstandalone_csrbank5_sel & builder_genericstandalone_interface5_bank_bus_we) & (builder_genericstandalone_interface5_bank_bus_adr[1:0] == 2'd2));
assign builder_genericstandalone_csrbank5_in_w = main_genericstandalone_i2c_status0[1:0];
assign main_genericstandalone_i2c_out_storage = main_genericstandalone_i2c_out_storage_full[1:0];
assign builder_genericstandalone_csrbank5_out0_w = main_genericstandalone_i2c_out_storage_full[1:0];
assign main_genericstandalone_i2c_oe_storage = main_genericstandalone_i2c_oe_storage_full[1:0];
assign builder_genericstandalone_csrbank5_oe0_w = main_genericstandalone_i2c_oe_storage_full[1:0];
assign builder_genericstandalone_csrbank6_sel = (builder_genericstandalone_interface6_bank_bus_adr[13:8] == 4'd10);
assign main_genericstandalone_genericstandalone_icap_iprog_r = builder_genericstandalone_interface6_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_icap_iprog_re = ((builder_genericstandalone_csrbank6_sel & builder_genericstandalone_interface6_bank_bus_we) & (builder_genericstandalone_interface6_bank_bus_adr[0] == 1'd0));
assign builder_genericstandalone_csrbank7_sel = (builder_genericstandalone_interface7_bank_bus_adr[13:8] == 2'd2);
assign builder_genericstandalone_csrbank7_address0_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_address0_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[0] == 1'd0));
assign builder_genericstandalone_csrbank7_data_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_data_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[0] == 1'd1));
assign main_genericstandalone_add_identifier_storage = main_genericstandalone_add_identifier_storage_full[7:0];
assign builder_genericstandalone_csrbank7_address0_w = main_genericstandalone_add_identifier_storage_full[7:0];
assign builder_genericstandalone_csrbank7_data_w = main_genericstandalone_add_identifier_status[7:0];
assign builder_genericstandalone_csrbank8_sel = (builder_genericstandalone_interface8_bank_bus_adr[13:8] == 4'd13);
assign builder_genericstandalone_csrbank8_reset0_r = builder_genericstandalone_interface8_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank8_reset0_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[0] == 1'd0));
assign main_genericstandalone_kernel_cpu_storage = main_genericstandalone_kernel_cpu_storage_full;
assign builder_genericstandalone_csrbank8_reset0_w = main_genericstandalone_kernel_cpu_storage_full;
assign builder_genericstandalone_csrbank9_sel = (builder_genericstandalone_interface9_bank_bus_adr[13:8] == 5'd18);
assign builder_genericstandalone_csrbank9_enable0_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank9_enable0_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 1'd0));
assign builder_genericstandalone_csrbank9_busy_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank9_busy_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 1'd1));
assign builder_genericstandalone_csrbank9_message_encoder_overflow_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank9_message_encoder_overflow_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 2'd2));
assign main_genericstandalone_rtio_analyzer_message_encoder_overflow_reset_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign main_genericstandalone_rtio_analyzer_message_encoder_overflow_reset_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 2'd3));
assign main_genericstandalone_rtio_analyzer_dma_reset_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign main_genericstandalone_rtio_analyzer_dma_reset_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 3'd4));
assign builder_genericstandalone_csrbank9_dma_base_address4_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank9_dma_base_address4_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 3'd5));
assign builder_genericstandalone_csrbank9_dma_base_address3_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_base_address3_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 3'd6));
assign builder_genericstandalone_csrbank9_dma_base_address2_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_base_address2_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 3'd7));
assign builder_genericstandalone_csrbank9_dma_base_address1_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_base_address1_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 4'd8));
assign builder_genericstandalone_csrbank9_dma_base_address0_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_base_address0_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 4'd9));
assign builder_genericstandalone_csrbank9_dma_last_address4_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank9_dma_last_address4_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 4'd10));
assign builder_genericstandalone_csrbank9_dma_last_address3_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_last_address3_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 4'd11));
assign builder_genericstandalone_csrbank9_dma_last_address2_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_last_address2_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 4'd12));
assign builder_genericstandalone_csrbank9_dma_last_address1_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_last_address1_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 4'd13));
assign builder_genericstandalone_csrbank9_dma_last_address0_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_last_address0_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 4'd14));
assign builder_genericstandalone_csrbank9_dma_byte_count7_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_byte_count7_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 4'd15));
assign builder_genericstandalone_csrbank9_dma_byte_count6_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_byte_count6_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 5'd16));
assign builder_genericstandalone_csrbank9_dma_byte_count5_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_byte_count5_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 5'd17));
assign builder_genericstandalone_csrbank9_dma_byte_count4_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_byte_count4_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 5'd18));
assign builder_genericstandalone_csrbank9_dma_byte_count3_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_byte_count3_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 5'd19));
assign builder_genericstandalone_csrbank9_dma_byte_count2_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_byte_count2_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 5'd20));
assign builder_genericstandalone_csrbank9_dma_byte_count1_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_byte_count1_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 5'd21));
assign builder_genericstandalone_csrbank9_dma_byte_count0_r = builder_genericstandalone_interface9_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank9_dma_byte_count0_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[4:0] == 5'd22));
assign main_genericstandalone_rtio_analyzer_enable_storage = main_genericstandalone_rtio_analyzer_enable_storage_full;
assign builder_genericstandalone_csrbank9_enable0_w = main_genericstandalone_rtio_analyzer_enable_storage_full;
assign builder_genericstandalone_csrbank9_busy_w = main_genericstandalone_rtio_analyzer_busy_status;
assign builder_genericstandalone_csrbank9_message_encoder_overflow_w = main_genericstandalone_rtio_analyzer_message_encoder_status;
assign main_genericstandalone_rtio_analyzer_dma_base_address_storage = main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[32:4];
assign builder_genericstandalone_csrbank9_dma_base_address4_w = main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[32];
assign builder_genericstandalone_csrbank9_dma_base_address3_w = main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[31:24];
assign builder_genericstandalone_csrbank9_dma_base_address2_w = main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[23:16];
assign builder_genericstandalone_csrbank9_dma_base_address1_w = main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[15:8];
assign builder_genericstandalone_csrbank9_dma_base_address0_w = {main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[7:4], {4{1'd0}}};
assign main_genericstandalone_rtio_analyzer_dma_last_address_storage = main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[32:4];
assign builder_genericstandalone_csrbank9_dma_last_address4_w = main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[32];
assign builder_genericstandalone_csrbank9_dma_last_address3_w = main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[31:24];
assign builder_genericstandalone_csrbank9_dma_last_address2_w = main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[23:16];
assign builder_genericstandalone_csrbank9_dma_last_address1_w = main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[15:8];
assign builder_genericstandalone_csrbank9_dma_last_address0_w = {main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[7:4], {4{1'd0}}};
assign builder_genericstandalone_csrbank9_dma_byte_count7_w = main_genericstandalone_rtio_analyzer_dma_status[63:56];
assign builder_genericstandalone_csrbank9_dma_byte_count6_w = main_genericstandalone_rtio_analyzer_dma_status[55:48];
assign builder_genericstandalone_csrbank9_dma_byte_count5_w = main_genericstandalone_rtio_analyzer_dma_status[47:40];
assign builder_genericstandalone_csrbank9_dma_byte_count4_w = main_genericstandalone_rtio_analyzer_dma_status[39:32];
assign builder_genericstandalone_csrbank9_dma_byte_count3_w = main_genericstandalone_rtio_analyzer_dma_status[31:24];
assign builder_genericstandalone_csrbank9_dma_byte_count2_w = main_genericstandalone_rtio_analyzer_dma_status[23:16];
assign builder_genericstandalone_csrbank9_dma_byte_count1_w = main_genericstandalone_rtio_analyzer_dma_status[15:8];
assign builder_genericstandalone_csrbank9_dma_byte_count0_w = main_genericstandalone_rtio_analyzer_dma_status[7:0];
assign builder_genericstandalone_csrbank10_sel = (builder_genericstandalone_interface10_bank_bus_adr[13:8] == 5'd16);
assign main_genericstandalone_rtio_core_reset_r = builder_genericstandalone_interface10_bank_bus_dat_w[0];
assign main_genericstandalone_rtio_core_reset_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 1'd0));
assign main_genericstandalone_rtio_core_reset_phy_r = builder_genericstandalone_interface10_bank_bus_dat_w[0];
assign main_genericstandalone_rtio_core_reset_phy_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 1'd1));
assign builder_genericstandalone_csrbank10_sed_spread_enable0_r = builder_genericstandalone_interface10_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank10_sed_spread_enable0_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 2'd2));
assign main_genericstandalone_rtio_core_async_error_r = builder_genericstandalone_interface10_bank_bus_dat_w[2:0];
assign main_genericstandalone_rtio_core_async_error_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 2'd3));
assign builder_genericstandalone_csrbank10_collision_channel1_r = builder_genericstandalone_interface10_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank10_collision_channel1_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 3'd4));
assign builder_genericstandalone_csrbank10_collision_channel0_r = builder_genericstandalone_interface10_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank10_collision_channel0_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 3'd5));
assign builder_genericstandalone_csrbank10_busy_channel1_r = builder_genericstandalone_interface10_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank10_busy_channel1_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 3'd6));
assign builder_genericstandalone_csrbank10_busy_channel0_r = builder_genericstandalone_interface10_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank10_busy_channel0_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 3'd7));
assign builder_genericstandalone_csrbank10_sequence_error_channel1_r = builder_genericstandalone_interface10_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank10_sequence_error_channel1_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 4'd8));
assign builder_genericstandalone_csrbank10_sequence_error_channel0_r = builder_genericstandalone_interface10_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank10_sequence_error_channel0_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[3:0] == 4'd9));
assign main_genericstandalone_rtio_core_storage = main_genericstandalone_rtio_core_storage_full;
assign builder_genericstandalone_csrbank10_sed_spread_enable0_w = main_genericstandalone_rtio_core_storage_full;
assign builder_genericstandalone_csrbank10_collision_channel1_w = main_genericstandalone_rtio_core_collision_channel_status[15:8];
assign builder_genericstandalone_csrbank10_collision_channel0_w = main_genericstandalone_rtio_core_collision_channel_status[7:0];
assign builder_genericstandalone_csrbank10_busy_channel1_w = main_genericstandalone_rtio_core_busy_channel_status[15:8];
assign builder_genericstandalone_csrbank10_busy_channel0_w = main_genericstandalone_rtio_core_busy_channel_status[7:0];
assign builder_genericstandalone_csrbank10_sequence_error_channel1_w = main_genericstandalone_rtio_core_sequence_error_channel_status[15:8];
assign builder_genericstandalone_csrbank10_sequence_error_channel0_w = main_genericstandalone_rtio_core_sequence_error_channel_status[7:0];
assign builder_genericstandalone_csrbank11_sel = (builder_genericstandalone_interface11_bank_bus_adr[13:8] == 5'd17);
assign builder_genericstandalone_csrbank11_mon_chan_sel0_r = builder_genericstandalone_interface11_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank11_mon_chan_sel0_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 1'd0));
assign builder_genericstandalone_csrbank11_mon_probe_sel0_r = builder_genericstandalone_interface11_bank_bus_dat_w[4:0];
assign builder_genericstandalone_csrbank11_mon_probe_sel0_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 1'd1));
assign main_genericstandalone_mon_value_update_r = builder_genericstandalone_interface11_bank_bus_dat_w[0];
assign main_genericstandalone_mon_value_update_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 2'd2));
assign builder_genericstandalone_csrbank11_mon_value3_r = builder_genericstandalone_interface11_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank11_mon_value3_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 2'd3));
assign builder_genericstandalone_csrbank11_mon_value2_r = builder_genericstandalone_interface11_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank11_mon_value2_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 3'd4));
assign builder_genericstandalone_csrbank11_mon_value1_r = builder_genericstandalone_interface11_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank11_mon_value1_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 3'd5));
assign builder_genericstandalone_csrbank11_mon_value0_r = builder_genericstandalone_interface11_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank11_mon_value0_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 3'd6));
assign builder_genericstandalone_csrbank11_inj_chan_sel0_r = builder_genericstandalone_interface11_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank11_inj_chan_sel0_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 3'd7));
assign builder_genericstandalone_csrbank11_inj_override_sel0_r = builder_genericstandalone_interface11_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank11_inj_override_sel0_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 4'd8));
assign main_genericstandalone_inj_value_r = builder_genericstandalone_interface11_bank_bus_dat_w[0];
assign main_genericstandalone_inj_value_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[3:0] == 4'd9));
assign main_genericstandalone_mon_chan_sel_storage = main_genericstandalone_mon_chan_sel_storage_full[5:0];
assign builder_genericstandalone_csrbank11_mon_chan_sel0_w = main_genericstandalone_mon_chan_sel_storage_full[5:0];
assign main_genericstandalone_mon_probe_sel_storage = main_genericstandalone_mon_probe_sel_storage_full[4:0];
assign builder_genericstandalone_csrbank11_mon_probe_sel0_w = main_genericstandalone_mon_probe_sel_storage_full[4:0];
assign builder_genericstandalone_csrbank11_mon_value3_w = main_genericstandalone_mon_status[31:24];
assign builder_genericstandalone_csrbank11_mon_value2_w = main_genericstandalone_mon_status[23:16];
assign builder_genericstandalone_csrbank11_mon_value1_w = main_genericstandalone_mon_status[15:8];
assign builder_genericstandalone_csrbank11_mon_value0_w = main_genericstandalone_mon_status[7:0];
assign main_genericstandalone_inj_chan_sel_storage = main_genericstandalone_inj_chan_sel_storage_full[5:0];
assign builder_genericstandalone_csrbank11_inj_chan_sel0_w = main_genericstandalone_inj_chan_sel_storage_full[5:0];
assign main_genericstandalone_inj_override_sel_storage = main_genericstandalone_inj_override_sel_storage_full[1:0];
assign builder_genericstandalone_csrbank11_inj_override_sel0_w = main_genericstandalone_inj_override_sel_storage_full[1:0];
assign builder_genericstandalone_csrbank12_sel = (builder_genericstandalone_interface12_bank_bus_adr[13:8] == 4'd9);
assign builder_genericstandalone_csrbank12_bitbang0_r = builder_genericstandalone_interface12_bank_bus_dat_w[3:0];
assign builder_genericstandalone_csrbank12_bitbang0_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[1:0] == 1'd0));
assign builder_genericstandalone_csrbank12_miso_r = builder_genericstandalone_interface12_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank12_miso_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[1:0] == 1'd1));
assign builder_genericstandalone_csrbank12_bitbang_en0_r = builder_genericstandalone_interface12_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank12_bitbang_en0_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[1:0] == 2'd2));
assign main_genericstandalone_genericstandalone_spiflash_bitbang_storage = main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full[3:0];
assign builder_genericstandalone_csrbank12_bitbang0_w = main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full[3:0];
assign builder_genericstandalone_csrbank12_miso_w = main_genericstandalone_genericstandalone_spiflash_status;
assign main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage = main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full;
assign builder_genericstandalone_csrbank12_bitbang_en0_w = main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full;
assign builder_genericstandalone_csrbank13_sel = (builder_genericstandalone_interface13_bank_bus_adr[13:8] == 2'd3);
assign builder_genericstandalone_csrbank13_load7_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_load7_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 1'd0));
assign builder_genericstandalone_csrbank13_load6_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_load6_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 1'd1));
assign builder_genericstandalone_csrbank13_load5_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_load5_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 2'd2));
assign builder_genericstandalone_csrbank13_load4_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_load4_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 2'd3));
assign builder_genericstandalone_csrbank13_load3_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_load3_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 3'd4));
assign builder_genericstandalone_csrbank13_load2_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_load2_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 3'd5));
assign builder_genericstandalone_csrbank13_load1_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_load1_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 3'd6));
assign builder_genericstandalone_csrbank13_load0_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_load0_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 3'd7));
assign builder_genericstandalone_csrbank13_reload7_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_reload7_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 4'd8));
assign builder_genericstandalone_csrbank13_reload6_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_reload6_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 4'd9));
assign builder_genericstandalone_csrbank13_reload5_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_reload5_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 4'd10));
assign builder_genericstandalone_csrbank13_reload4_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_reload4_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 4'd11));
assign builder_genericstandalone_csrbank13_reload3_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_reload3_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 4'd12));
assign builder_genericstandalone_csrbank13_reload2_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_reload2_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 4'd13));
assign builder_genericstandalone_csrbank13_reload1_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_reload1_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 4'd14));
assign builder_genericstandalone_csrbank13_reload0_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_reload0_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 4'd15));
assign builder_genericstandalone_csrbank13_en0_r = builder_genericstandalone_interface13_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank13_en0_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd16));
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_r = builder_genericstandalone_interface13_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd17));
assign builder_genericstandalone_csrbank13_value7_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_value7_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd18));
assign builder_genericstandalone_csrbank13_value6_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_value6_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd19));
assign builder_genericstandalone_csrbank13_value5_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_value5_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd20));
assign builder_genericstandalone_csrbank13_value4_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_value4_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd21));
assign builder_genericstandalone_csrbank13_value3_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_value3_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd22));
assign builder_genericstandalone_csrbank13_value2_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_value2_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd23));
assign builder_genericstandalone_csrbank13_value1_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_value1_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd24));
assign builder_genericstandalone_csrbank13_value0_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_value0_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd25));
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_r = builder_genericstandalone_interface13_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd26));
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_r = builder_genericstandalone_interface13_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd27));
assign builder_genericstandalone_csrbank13_ev_enable0_r = builder_genericstandalone_interface13_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank13_ev_enable0_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[4:0] == 5'd28));
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[63:0];
assign builder_genericstandalone_csrbank13_load7_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[63:56];
assign builder_genericstandalone_csrbank13_load6_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[55:48];
assign builder_genericstandalone_csrbank13_load5_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[47:40];
assign builder_genericstandalone_csrbank13_load4_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[39:32];
assign builder_genericstandalone_csrbank13_load3_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[31:24];
assign builder_genericstandalone_csrbank13_load2_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[23:16];
assign builder_genericstandalone_csrbank13_load1_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[15:8];
assign builder_genericstandalone_csrbank13_load0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[63:0];
assign builder_genericstandalone_csrbank13_reload7_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[63:56];
assign builder_genericstandalone_csrbank13_reload6_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[55:48];
assign builder_genericstandalone_csrbank13_reload5_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[47:40];
assign builder_genericstandalone_csrbank13_reload4_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[39:32];
assign builder_genericstandalone_csrbank13_reload3_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[31:24];
assign builder_genericstandalone_csrbank13_reload2_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[23:16];
assign builder_genericstandalone_csrbank13_reload1_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[15:8];
assign builder_genericstandalone_csrbank13_reload0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage = main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full;
assign builder_genericstandalone_csrbank13_en0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full;
assign builder_genericstandalone_csrbank13_value7_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[63:56];
assign builder_genericstandalone_csrbank13_value6_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[55:48];
assign builder_genericstandalone_csrbank13_value5_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[47:40];
assign builder_genericstandalone_csrbank13_value4_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[39:32];
assign builder_genericstandalone_csrbank13_value3_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[31:24];
assign builder_genericstandalone_csrbank13_value2_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[23:16];
assign builder_genericstandalone_csrbank13_value1_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[15:8];
assign builder_genericstandalone_csrbank13_value0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage = main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full;
assign builder_genericstandalone_csrbank13_ev_enable0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full;
assign builder_genericstandalone_csrbank14_sel = (builder_genericstandalone_interface14_bank_bus_adr[13:8] == 1'd1);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_r = builder_genericstandalone_interface14_bank_bus_dat_w[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 1'd0));
assign builder_genericstandalone_csrbank14_txfull_r = builder_genericstandalone_interface14_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank14_txfull_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 1'd1));
assign builder_genericstandalone_csrbank14_rxempty_r = builder_genericstandalone_interface14_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank14_rxempty_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 2'd2));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_status_r = builder_genericstandalone_interface14_bank_bus_dat_w[1:0];
assign main_genericstandalone_genericstandalone_genericstandalone_uart_status_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 2'd3));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_pending_r = builder_genericstandalone_interface14_bank_bus_dat_w[1:0];
assign main_genericstandalone_genericstandalone_genericstandalone_uart_pending_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 3'd4));
assign builder_genericstandalone_csrbank14_ev_enable0_r = builder_genericstandalone_interface14_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank14_ev_enable0_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 3'd5));
assign builder_genericstandalone_csrbank14_txfull_w = main_genericstandalone_genericstandalone_genericstandalone_uart_txfull_status;
assign builder_genericstandalone_csrbank14_rxempty_w = main_genericstandalone_genericstandalone_genericstandalone_uart_rxempty_status;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_storage = main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full[1:0];
assign builder_genericstandalone_csrbank14_ev_enable0_w = main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full[1:0];
assign builder_genericstandalone_csrbank15_sel = (builder_genericstandalone_interface15_bank_bus_adr[13:8] == 1'd0);
assign builder_genericstandalone_csrbank15_tuning_word3_r = builder_genericstandalone_interface15_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank15_tuning_word3_re = ((builder_genericstandalone_csrbank15_sel & builder_genericstandalone_interface15_bank_bus_we) & (builder_genericstandalone_interface15_bank_bus_adr[1:0] == 1'd0));
assign builder_genericstandalone_csrbank15_tuning_word2_r = builder_genericstandalone_interface15_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank15_tuning_word2_re = ((builder_genericstandalone_csrbank15_sel & builder_genericstandalone_interface15_bank_bus_we) & (builder_genericstandalone_interface15_bank_bus_adr[1:0] == 1'd1));
assign builder_genericstandalone_csrbank15_tuning_word1_r = builder_genericstandalone_interface15_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank15_tuning_word1_re = ((builder_genericstandalone_csrbank15_sel & builder_genericstandalone_interface15_bank_bus_we) & (builder_genericstandalone_interface15_bank_bus_adr[1:0] == 2'd2));
assign builder_genericstandalone_csrbank15_tuning_word0_r = builder_genericstandalone_interface15_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank15_tuning_word0_re = ((builder_genericstandalone_csrbank15_sel & builder_genericstandalone_interface15_bank_bus_we) & (builder_genericstandalone_interface15_bank_bus_adr[1:0] == 2'd3));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[31:0];
assign builder_genericstandalone_csrbank15_tuning_word3_w = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[31:24];
assign builder_genericstandalone_csrbank15_tuning_word2_w = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[23:16];
assign builder_genericstandalone_csrbank15_tuning_word1_w = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[15:8];
assign builder_genericstandalone_csrbank15_tuning_word0_w = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[7:0];
assign builder_genericstandalone_csrbank16_sel = (builder_genericstandalone_interface16_bank_bus_adr[13:8] == 4'd8);
assign builder_genericstandalone_csrbank16_status_r = builder_genericstandalone_interface16_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank16_status_re = ((builder_genericstandalone_csrbank16_sel & builder_genericstandalone_interface16_bank_bus_we) & (builder_genericstandalone_interface16_bank_bus_adr[0] == 1'd0));
assign builder_genericstandalone_csrbank16_status_w = main_genericstandalone_genericstandalone_virtual_leds_status[7:0];
assign builder_genericstandalone_interface0_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface1_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface2_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface3_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface4_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface5_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface6_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface7_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface8_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface9_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface10_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface11_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface12_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface13_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface14_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface15_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface16_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface0_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface1_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface2_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface3_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface4_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface5_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface6_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface7_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface8_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface9_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface10_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface11_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface12_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface13_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface14_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface15_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface16_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface0_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface1_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface2_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface3_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface4_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface5_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface6_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface7_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface8_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface9_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface10_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface11_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface12_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface13_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface14_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface15_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface16_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_interface_dat_r = ((((((((((((((((builder_genericstandalone_interface0_bank_bus_dat_r | builder_genericstandalone_interface1_bank_bus_dat_r) | builder_genericstandalone_interface2_bank_bus_dat_r) | builder_genericstandalone_interface3_bank_bus_dat_r) | builder_genericstandalone_interface4_bank_bus_dat_r) | builder_genericstandalone_interface5_bank_bus_dat_r) | builder_genericstandalone_interface6_bank_bus_dat_r) | builder_genericstandalone_interface7_bank_bus_dat_r) | builder_genericstandalone_interface8_bank_bus_dat_r) | builder_genericstandalone_interface9_bank_bus_dat_r) | builder_genericstandalone_interface10_bank_bus_dat_r) | builder_genericstandalone_interface11_bank_bus_dat_r) | builder_genericstandalone_interface12_bank_bus_dat_r) | builder_genericstandalone_interface13_bank_bus_dat_r) | builder_genericstandalone_interface14_bank_bus_dat_r) | builder_genericstandalone_interface15_bank_bus_dat_r) | builder_genericstandalone_interface16_bank_bus_dat_r);
assign builder_slice_proxy0 = main_genericstandalone_interface0_bus_dat_r[63:0];
assign builder_slice_proxy1 = main_genericstandalone_interface0_bus_dat_r[63:0];
assign builder_slice_proxy2 = main_genericstandalone_interface0_bus_dat_r[63:0];
assign builder_slice_proxy3 = main_genericstandalone_interface0_bus_dat_r[63:0];
assign builder_slice_proxy4 = main_genericstandalone_interface0_bus_dat_r[63:0];
assign builder_slice_proxy5 = main_genericstandalone_interface0_bus_dat_r[63:0];
assign builder_slice_proxy6 = main_genericstandalone_interface0_bus_dat_r[63:0];
assign builder_slice_proxy7 = main_genericstandalone_interface0_bus_dat_r[63:0];
assign builder_slice_proxy8 = main_genericstandalone_interface0_bus_dat_r[127:64];
assign builder_slice_proxy9 = main_genericstandalone_interface0_bus_dat_r[127:64];
assign builder_slice_proxy10 = main_genericstandalone_interface0_bus_dat_r[127:64];
assign builder_slice_proxy11 = main_genericstandalone_interface0_bus_dat_r[127:64];
assign builder_slice_proxy12 = main_genericstandalone_interface0_bus_dat_r[127:64];
assign builder_slice_proxy13 = main_genericstandalone_interface0_bus_dat_r[127:64];
assign builder_slice_proxy14 = main_genericstandalone_interface0_bus_dat_r[127:64];
assign builder_slice_proxy15 = main_genericstandalone_interface0_bus_dat_r[127:64];
assign builder_slice_proxy16 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[63:0];
assign builder_slice_proxy17 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[63:0];
assign builder_slice_proxy18 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[63:0];
assign builder_slice_proxy19 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[63:0];
assign builder_slice_proxy20 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[63:0];
assign builder_slice_proxy21 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[63:0];
assign builder_slice_proxy22 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[63:0];
assign builder_slice_proxy23 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[63:0];
assign builder_slice_proxy24 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[127:64];
assign builder_slice_proxy25 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[127:64];
assign builder_slice_proxy26 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[127:64];
assign builder_slice_proxy27 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[127:64];
assign builder_slice_proxy28 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[127:64];
assign builder_slice_proxy29 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[127:64];
assign builder_slice_proxy30 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[127:64];
assign builder_slice_proxy31 = main_genericstandalone_rtio_analyzer_dma_sink_payload_data[127:64];

// synthesis translate_off
reg dummy_d_221;
// synthesis translate_on
always @(*) begin
	builder_comb_basiclowerer_self <= 32'd0;
	case (main_genericstandalone_genericstandalone_icap_counter1)
		1'd0: begin
			builder_comb_basiclowerer_self <= 32'd4294967295;
		end
		1'd1: begin
			builder_comb_basiclowerer_self <= 8'd187;
		end
		2'd2: begin
			builder_comb_basiclowerer_self <= 29'd287440964;
		end
		2'd3: begin
			builder_comb_basiclowerer_self <= 32'd4294967295;
		end
		3'd4: begin
			builder_comb_basiclowerer_self <= 31'd1436133990;
		end
		3'd5: begin
			builder_comb_basiclowerer_self <= 27'd67108864;
		end
		3'd6: begin
			builder_comb_basiclowerer_self <= 28'd205521024;
		end
		3'd7: begin
			builder_comb_basiclowerer_self <= 1'd0;
		end
		4'd8: begin
			builder_comb_basiclowerer_self <= 28'd201326976;
		end
		4'd9: begin
			builder_comb_basiclowerer_self <= 8'd240;
		end
		default: begin
			builder_comb_basiclowerer_self <= 27'd67108864;
		end
	endcase
// synthesis translate_off
	dummy_d_221 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_222;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self0 <= 29'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_self0 <= main_genericstandalone_kernel_cpu_ibus_adr;
		end
		default: begin
			builder_comb_rhs_self0 <= main_genericstandalone_kernel_cpu_dbus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_222 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_223;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self1 <= 64'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_self1 <= main_genericstandalone_kernel_cpu_ibus_dat_w;
		end
		default: begin
			builder_comb_rhs_self1 <= main_genericstandalone_kernel_cpu_dbus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_223 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_224;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self2 <= 8'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_self2 <= main_genericstandalone_kernel_cpu_ibus_sel;
		end
		default: begin
			builder_comb_rhs_self2 <= main_genericstandalone_kernel_cpu_dbus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_224 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_225;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self3 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_self3 <= main_genericstandalone_kernel_cpu_ibus_cyc;
		end
		default: begin
			builder_comb_rhs_self3 <= main_genericstandalone_kernel_cpu_dbus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_225 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_226;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self4 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_self4 <= main_genericstandalone_kernel_cpu_ibus_stb;
		end
		default: begin
			builder_comb_rhs_self4 <= main_genericstandalone_kernel_cpu_dbus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_226 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_227;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self5 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_self5 <= main_genericstandalone_kernel_cpu_ibus_we;
		end
		default: begin
			builder_comb_rhs_self5 <= main_genericstandalone_kernel_cpu_dbus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_227 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_228;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self6 <= 3'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_self6 <= main_genericstandalone_kernel_cpu_ibus_cti;
		end
		default: begin
			builder_comb_rhs_self6 <= main_genericstandalone_kernel_cpu_dbus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_228 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_229;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self7 <= 2'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_self7 <= main_genericstandalone_kernel_cpu_ibus_bte;
		end
		default: begin
			builder_comb_rhs_self7 <= main_genericstandalone_kernel_cpu_dbus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_229 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_230;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self8 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_lane_dist_current_lane)
		1'd0: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record0_high_watermark;
		end
		1'd1: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record1_high_watermark;
		end
		2'd2: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record2_high_watermark;
		end
		2'd3: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record3_high_watermark;
		end
		3'd4: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record4_high_watermark;
		end
		3'd5: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record5_high_watermark;
		end
		3'd6: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record6_high_watermark;
		end
		3'd7: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record7_high_watermark;
		end
		4'd8: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record8_high_watermark;
		end
		4'd9: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record9_high_watermark;
		end
		4'd10: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record10_high_watermark;
		end
		4'd11: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record11_high_watermark;
		end
		4'd12: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record12_high_watermark;
		end
		4'd13: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record13_high_watermark;
		end
		4'd14: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record14_high_watermark;
		end
		default: begin
			builder_comb_rhs_self8 <= main_genericstandalone_rtio_core_sed_lane_dist_record15_high_watermark;
		end
	endcase
// synthesis translate_off
	dummy_d_230 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_231;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self9 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_lane_dist_current_lane)
		1'd0: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record0_writable;
		end
		1'd1: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record1_writable;
		end
		2'd2: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record2_writable;
		end
		2'd3: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record3_writable;
		end
		3'd4: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record4_writable;
		end
		3'd5: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record5_writable;
		end
		3'd6: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record6_writable;
		end
		3'd7: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record7_writable;
		end
		4'd8: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record8_writable;
		end
		4'd9: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record9_writable;
		end
		4'd10: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record10_writable;
		end
		4'd11: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record11_writable;
		end
		4'd12: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record12_writable;
		end
		4'd13: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record13_writable;
		end
		4'd14: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record14_writable;
		end
		default: begin
			builder_comb_rhs_self9 <= main_genericstandalone_rtio_core_sed_lane_dist_record15_writable;
		end
	endcase
// synthesis translate_off
	dummy_d_231 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_232;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self10 <= 2'd0;
	case (main_genericstandalone_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow0, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow0))};
		end
		1'd1: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow1, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow1))};
		end
		2'd2: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow2, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow2))};
		end
		2'd3: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow3, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow3))};
		end
		3'd4: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		3'd5: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		3'd6: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		3'd7: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		4'd8: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		4'd9: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		4'd10: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		4'd11: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		4'd12: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		4'd13: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		4'd14: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		4'd15: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd16: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow4, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow4))};
		end
		5'd17: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd18: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd19: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd20: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd21: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd22: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow5, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow5))};
		end
		5'd23: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd24: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd25: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd26: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd27: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd28: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow6, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow6))};
		end
		5'd29: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow7, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow7))};
		end
		5'd30: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		5'd31: begin
			builder_comb_rhs_self10 <= {main_genericstandalone_rtio_core_inputcollector_overflow8, (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_readable & (~main_genericstandalone_rtio_core_inputcollector_overflow8))};
		end
		6'd32: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		6'd33: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		6'd34: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		6'd35: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		6'd36: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_self10 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_232 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_233;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self11 <= 2'd0;
	case (main_genericstandalone_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_self11 <= main_genericstandalone_rtio_cri_cmd;
		end
		default: begin
			builder_comb_rhs_self11 <= main_genericstandalone_dma_cri_master_cri_cmd;
		end
	endcase
// synthesis translate_off
	dummy_d_233 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_234;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self12 <= 24'd0;
	case (main_genericstandalone_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_self12 <= main_genericstandalone_rtio_cri_chan_sel;
		end
		default: begin
			builder_comb_rhs_self12 <= main_genericstandalone_dma_cri_master_cri_chan_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_234 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_235;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self13 <= 64'd0;
	case (main_genericstandalone_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_self13 <= main_genericstandalone_rtio_cri_o_timestamp;
		end
		default: begin
			builder_comb_rhs_self13 <= main_genericstandalone_dma_cri_master_cri_o_timestamp;
		end
	endcase
// synthesis translate_off
	dummy_d_235 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_236;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self14 <= 512'd0;
	case (main_genericstandalone_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_self14 <= main_genericstandalone_rtio_cri_o_data;
		end
		default: begin
			builder_comb_rhs_self14 <= main_genericstandalone_dma_cri_master_cri_o_data;
		end
	endcase
// synthesis translate_off
	dummy_d_236 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_237;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self15 <= 8'd0;
	case (main_genericstandalone_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_self15 <= main_genericstandalone_rtio_cri_o_address;
		end
		default: begin
			builder_comb_rhs_self15 <= main_genericstandalone_dma_cri_master_cri_o_address;
		end
	endcase
// synthesis translate_off
	dummy_d_237 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_238;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self16 <= 64'd0;
	case (main_genericstandalone_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_self16 <= main_genericstandalone_rtio_cri_i_timeout;
		end
		default: begin
			builder_comb_rhs_self16 <= main_genericstandalone_dma_cri_master_cri_i_timeout;
		end
	endcase
// synthesis translate_off
	dummy_d_238 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_239;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self18 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self18 <= main_genericstandalone_inj_o_sys0;
		end
		1'd1: begin
			builder_comb_rhs_self18 <= main_genericstandalone_inj_o_sys1;
		end
		default: begin
			builder_comb_rhs_self18 <= main_genericstandalone_inj_o_sys2;
		end
	endcase
// synthesis translate_off
	dummy_d_239 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_240;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self19 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self19 <= main_genericstandalone_inj_o_sys3;
		end
		1'd1: begin
			builder_comb_rhs_self19 <= main_genericstandalone_inj_o_sys4;
		end
		default: begin
			builder_comb_rhs_self19 <= main_genericstandalone_inj_o_sys5;
		end
	endcase
// synthesis translate_off
	dummy_d_240 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_241;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self20 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self20 <= main_genericstandalone_inj_o_sys6;
		end
		1'd1: begin
			builder_comb_rhs_self20 <= main_genericstandalone_inj_o_sys7;
		end
		default: begin
			builder_comb_rhs_self20 <= main_genericstandalone_inj_o_sys8;
		end
	endcase
// synthesis translate_off
	dummy_d_241 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_242;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self21 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self21 <= main_genericstandalone_inj_o_sys9;
		end
		1'd1: begin
			builder_comb_rhs_self21 <= main_genericstandalone_inj_o_sys10;
		end
		default: begin
			builder_comb_rhs_self21 <= main_genericstandalone_inj_o_sys11;
		end
	endcase
// synthesis translate_off
	dummy_d_242 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_243;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self22 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self22 <= main_genericstandalone_inj_o_sys12;
		end
		1'd1: begin
			builder_comb_rhs_self22 <= main_genericstandalone_inj_o_sys13;
		end
		default: begin
			builder_comb_rhs_self22 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_243 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_244;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self23 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self23 <= main_genericstandalone_inj_o_sys14;
		end
		1'd1: begin
			builder_comb_rhs_self23 <= main_genericstandalone_inj_o_sys15;
		end
		default: begin
			builder_comb_rhs_self23 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_244 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_245;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self24 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self24 <= main_genericstandalone_inj_o_sys16;
		end
		1'd1: begin
			builder_comb_rhs_self24 <= main_genericstandalone_inj_o_sys17;
		end
		default: begin
			builder_comb_rhs_self24 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_245 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_246;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self25 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self25 <= main_genericstandalone_inj_o_sys18;
		end
		1'd1: begin
			builder_comb_rhs_self25 <= main_genericstandalone_inj_o_sys19;
		end
		default: begin
			builder_comb_rhs_self25 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_246 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_247;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self26 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self26 <= main_genericstandalone_inj_o_sys20;
		end
		1'd1: begin
			builder_comb_rhs_self26 <= main_genericstandalone_inj_o_sys21;
		end
		default: begin
			builder_comb_rhs_self26 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_247 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_248;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self27 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self27 <= main_genericstandalone_inj_o_sys22;
		end
		1'd1: begin
			builder_comb_rhs_self27 <= main_genericstandalone_inj_o_sys23;
		end
		default: begin
			builder_comb_rhs_self27 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_248 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_249;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self28 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self28 <= main_genericstandalone_inj_o_sys24;
		end
		1'd1: begin
			builder_comb_rhs_self28 <= main_genericstandalone_inj_o_sys25;
		end
		default: begin
			builder_comb_rhs_self28 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_249 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_250;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self29 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self29 <= main_genericstandalone_inj_o_sys26;
		end
		1'd1: begin
			builder_comb_rhs_self29 <= main_genericstandalone_inj_o_sys27;
		end
		default: begin
			builder_comb_rhs_self29 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_250 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_251;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self30 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self30 <= main_genericstandalone_inj_o_sys28;
		end
		1'd1: begin
			builder_comb_rhs_self30 <= main_genericstandalone_inj_o_sys29;
		end
		default: begin
			builder_comb_rhs_self30 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_251 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_252;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self31 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self31 <= main_genericstandalone_inj_o_sys30;
		end
		1'd1: begin
			builder_comb_rhs_self31 <= main_genericstandalone_inj_o_sys31;
		end
		default: begin
			builder_comb_rhs_self31 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_252 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_253;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self32 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self32 <= main_genericstandalone_inj_o_sys32;
		end
		1'd1: begin
			builder_comb_rhs_self32 <= main_genericstandalone_inj_o_sys33;
		end
		default: begin
			builder_comb_rhs_self32 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_253 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_254;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self33 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self33 <= main_genericstandalone_inj_o_sys34;
		end
		1'd1: begin
			builder_comb_rhs_self33 <= main_genericstandalone_inj_o_sys35;
		end
		default: begin
			builder_comb_rhs_self33 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_254 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_255;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self34 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self34 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_self34 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_self34 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_255 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_256;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self35 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self35 <= main_genericstandalone_inj_o_sys36;
		end
		1'd1: begin
			builder_comb_rhs_self35 <= main_genericstandalone_inj_o_sys37;
		end
		default: begin
			builder_comb_rhs_self35 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_256 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_257;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self36 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self36 <= main_genericstandalone_inj_o_sys38;
		end
		1'd1: begin
			builder_comb_rhs_self36 <= main_genericstandalone_inj_o_sys39;
		end
		default: begin
			builder_comb_rhs_self36 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_257 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_258;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self37 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self37 <= main_genericstandalone_inj_o_sys40;
		end
		1'd1: begin
			builder_comb_rhs_self37 <= main_genericstandalone_inj_o_sys41;
		end
		default: begin
			builder_comb_rhs_self37 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_258 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_259;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self38 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self38 <= main_genericstandalone_inj_o_sys42;
		end
		1'd1: begin
			builder_comb_rhs_self38 <= main_genericstandalone_inj_o_sys43;
		end
		default: begin
			builder_comb_rhs_self38 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_259 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_260;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self39 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self39 <= main_genericstandalone_inj_o_sys44;
		end
		1'd1: begin
			builder_comb_rhs_self39 <= main_genericstandalone_inj_o_sys45;
		end
		default: begin
			builder_comb_rhs_self39 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_260 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_261;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self40 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self40 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_self40 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_self40 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_261 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_262;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self41 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self41 <= main_genericstandalone_inj_o_sys46;
		end
		1'd1: begin
			builder_comb_rhs_self41 <= main_genericstandalone_inj_o_sys47;
		end
		default: begin
			builder_comb_rhs_self41 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_262 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_263;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self42 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self42 <= main_genericstandalone_inj_o_sys48;
		end
		1'd1: begin
			builder_comb_rhs_self42 <= main_genericstandalone_inj_o_sys49;
		end
		default: begin
			builder_comb_rhs_self42 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_263 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_264;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self43 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self43 <= main_genericstandalone_inj_o_sys50;
		end
		1'd1: begin
			builder_comb_rhs_self43 <= main_genericstandalone_inj_o_sys51;
		end
		default: begin
			builder_comb_rhs_self43 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_264 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_265;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self44 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self44 <= main_genericstandalone_inj_o_sys52;
		end
		1'd1: begin
			builder_comb_rhs_self44 <= main_genericstandalone_inj_o_sys53;
		end
		default: begin
			builder_comb_rhs_self44 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_265 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_266;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self45 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self45 <= main_genericstandalone_inj_o_sys54;
		end
		1'd1: begin
			builder_comb_rhs_self45 <= main_genericstandalone_inj_o_sys55;
		end
		default: begin
			builder_comb_rhs_self45 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_266 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_267;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self46 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self46 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_self46 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_self46 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_267 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_268;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self47 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self47 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_self47 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_self47 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_268 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_269;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self48 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self48 <= main_genericstandalone_inj_o_sys56;
		end
		1'd1: begin
			builder_comb_rhs_self48 <= main_genericstandalone_inj_o_sys57;
		end
		default: begin
			builder_comb_rhs_self48 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_269 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_270;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self49 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self49 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_self49 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_self49 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_270 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_271;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self50 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self50 <= main_genericstandalone_inj_o_sys58;
		end
		1'd1: begin
			builder_comb_rhs_self50 <= main_genericstandalone_inj_o_sys59;
		end
		default: begin
			builder_comb_rhs_self50 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_271 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_272;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self51 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self51 <= main_genericstandalone_inj_o_sys60;
		end
		1'd1: begin
			builder_comb_rhs_self51 <= main_genericstandalone_inj_o_sys61;
		end
		default: begin
			builder_comb_rhs_self51 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_272 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_273;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self52 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self52 <= main_genericstandalone_inj_o_sys62;
		end
		1'd1: begin
			builder_comb_rhs_self52 <= main_genericstandalone_inj_o_sys63;
		end
		default: begin
			builder_comb_rhs_self52 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_273 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_274;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self53 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self53 <= main_genericstandalone_inj_o_sys64;
		end
		1'd1: begin
			builder_comb_rhs_self53 <= main_genericstandalone_inj_o_sys65;
		end
		default: begin
			builder_comb_rhs_self53 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_274 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_275;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self54 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self54 <= main_genericstandalone_inj_o_sys66;
		end
		1'd1: begin
			builder_comb_rhs_self54 <= main_genericstandalone_inj_o_sys67;
		end
		default: begin
			builder_comb_rhs_self54 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_275 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_276;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self55 <= 1'd0;
	case (main_genericstandalone_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_self55 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_self55 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_self55 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_276 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_277;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self17 <= 1'd0;
	case (main_genericstandalone_inj_chan_sel_storage)
		1'd0: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self18;
		end
		1'd1: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self19;
		end
		2'd2: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self20;
		end
		2'd3: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self21;
		end
		3'd4: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self22;
		end
		3'd5: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self23;
		end
		3'd6: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self24;
		end
		3'd7: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self25;
		end
		4'd8: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self26;
		end
		4'd9: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self27;
		end
		4'd10: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self28;
		end
		4'd11: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self29;
		end
		4'd12: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self30;
		end
		4'd13: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self31;
		end
		4'd14: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self32;
		end
		4'd15: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self33;
		end
		5'd16: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self34;
		end
		5'd17: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self35;
		end
		5'd18: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self36;
		end
		5'd19: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self37;
		end
		5'd20: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self38;
		end
		5'd21: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self39;
		end
		5'd22: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self40;
		end
		5'd23: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self41;
		end
		5'd24: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self42;
		end
		5'd25: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self43;
		end
		5'd26: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self44;
		end
		5'd27: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self45;
		end
		5'd28: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self46;
		end
		5'd29: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self47;
		end
		5'd30: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self48;
		end
		5'd31: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self49;
		end
		6'd32: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self50;
		end
		6'd33: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self51;
		end
		6'd34: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self52;
		end
		6'd35: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self53;
		end
		6'd36: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self54;
		end
		default: begin
			builder_comb_rhs_self17 <= builder_comb_rhs_self55;
		end
	endcase
// synthesis translate_off
	dummy_d_277 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_278;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self56 <= 29'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self56 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_adr;
		end
		default: begin
			builder_comb_rhs_self56 <= main_genericstandalone_kernel_cpu_wb_sdram_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_278 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_279;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self57 <= 64'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self57 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_w;
		end
		default: begin
			builder_comb_rhs_self57 <= main_genericstandalone_kernel_cpu_wb_sdram_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_279 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_280;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self58 <= 8'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self58 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_sel;
		end
		default: begin
			builder_comb_rhs_self58 <= main_genericstandalone_kernel_cpu_wb_sdram_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_280 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_281;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self59 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self59 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cyc;
		end
		default: begin
			builder_comb_rhs_self59 <= main_genericstandalone_kernel_cpu_wb_sdram_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_281 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_282;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self60 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self60 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_stb;
		end
		default: begin
			builder_comb_rhs_self60 <= main_genericstandalone_kernel_cpu_wb_sdram_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_282 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_283;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self61 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self61 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_we;
		end
		default: begin
			builder_comb_rhs_self61 <= main_genericstandalone_kernel_cpu_wb_sdram_we;
		end
	endcase
// synthesis translate_off
	dummy_d_283 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_284;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self62 <= 3'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self62 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cti;
		end
		default: begin
			builder_comb_rhs_self62 <= main_genericstandalone_kernel_cpu_wb_sdram_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_284 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_285;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self63 <= 2'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self63 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_bte;
		end
		default: begin
			builder_comb_rhs_self63 <= main_genericstandalone_kernel_cpu_wb_sdram_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_285 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_286;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self64 <= 29'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self64 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_adr;
		end
		1'd1: begin
			builder_comb_rhs_self64 <= main_genericstandalone_interface0_bus_adr;
		end
		default: begin
			builder_comb_rhs_self64 <= main_genericstandalone_interface1_bus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_286 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_287;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self65 <= 128'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self65 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w;
		end
		1'd1: begin
			builder_comb_rhs_self65 <= main_genericstandalone_interface0_bus_dat_w;
		end
		default: begin
			builder_comb_rhs_self65 <= main_genericstandalone_interface1_bus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_287 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_288;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self66 <= 16'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self66 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_sel;
		end
		1'd1: begin
			builder_comb_rhs_self66 <= main_genericstandalone_interface0_bus_sel;
		end
		default: begin
			builder_comb_rhs_self66 <= main_genericstandalone_interface1_bus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_288 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_289;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self67 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self67 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc;
		end
		1'd1: begin
			builder_comb_rhs_self67 <= main_genericstandalone_interface0_bus_cyc;
		end
		default: begin
			builder_comb_rhs_self67 <= main_genericstandalone_interface1_bus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_289 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_290;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self68 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self68 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb;
		end
		1'd1: begin
			builder_comb_rhs_self68 <= main_genericstandalone_interface0_bus_stb;
		end
		default: begin
			builder_comb_rhs_self68 <= main_genericstandalone_interface1_bus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_290 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_291;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self69 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self69 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we;
		end
		1'd1: begin
			builder_comb_rhs_self69 <= main_genericstandalone_interface0_bus_we;
		end
		default: begin
			builder_comb_rhs_self69 <= main_genericstandalone_interface1_bus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_291 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_292;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self70 <= 3'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self70 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cti;
		end
		1'd1: begin
			builder_comb_rhs_self70 <= main_genericstandalone_interface0_bus_cti;
		end
		default: begin
			builder_comb_rhs_self70 <= main_genericstandalone_interface1_bus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_292 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_293;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self71 <= 2'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_self71 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_bte;
		end
		1'd1: begin
			builder_comb_rhs_self71 <= main_genericstandalone_interface0_bus_bte;
		end
		default: begin
			builder_comb_rhs_self71 <= main_genericstandalone_interface1_bus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_293 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_294;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self72 <= 29'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_self72 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_adr;
		end
		default: begin
			builder_comb_rhs_self72 <= main_genericstandalone_genericstandalone_genericstandalone_dbus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_294 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_295;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self73 <= 64'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_self73 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_w;
		end
		default: begin
			builder_comb_rhs_self73 <= main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_295 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_296;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self74 <= 8'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_self74 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_sel;
		end
		default: begin
			builder_comb_rhs_self74 <= main_genericstandalone_genericstandalone_genericstandalone_dbus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_296 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_297;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self75 <= 1'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_self75 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_cyc;
		end
		default: begin
			builder_comb_rhs_self75 <= main_genericstandalone_genericstandalone_genericstandalone_dbus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_297 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_298;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self76 <= 1'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_self76 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_stb;
		end
		default: begin
			builder_comb_rhs_self76 <= main_genericstandalone_genericstandalone_genericstandalone_dbus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_298 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_299;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self77 <= 1'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_self77 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_we;
		end
		default: begin
			builder_comb_rhs_self77 <= main_genericstandalone_genericstandalone_genericstandalone_dbus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_299 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_300;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self78 <= 3'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_self78 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_cti;
		end
		default: begin
			builder_comb_rhs_self78 <= main_genericstandalone_genericstandalone_genericstandalone_dbus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_300 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_301;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_self79 <= 2'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_self79 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_bte;
		end
		default: begin
			builder_comb_rhs_self79 <= main_genericstandalone_genericstandalone_genericstandalone_dbus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_301 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_302;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self0 <= 3'd0;
	case (main_genericstandalone_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self0 <= 3'd4;
		end
		2'd3: begin
			builder_sync_t_rhs_self0 <= 2'd3;
		end
		3'd4: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self0 <= 2'd2;
		end
		3'd6: begin
			builder_sync_t_rhs_self0 <= 3'd6;
		end
		3'd7: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self0 <= 3'd7;
		end
		4'd9: begin
			builder_sync_t_rhs_self0 <= 1'd1;
		end
		4'd10: begin
			builder_sync_t_rhs_self0 <= 3'd5;
		end
		4'd11: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_302 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_303;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self0 <= 3'd0;
	case (main_genericstandalone_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
		2'd2: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
		2'd3: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
		3'd4: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_f_t_self0 <= 3'd5;
		end
		3'd6: begin
			builder_sync_f_t_self0 <= 1'd1;
		end
		3'd7: begin
			builder_sync_f_t_self0 <= 3'd7;
		end
		4'd8: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
		4'd9: begin
			builder_sync_f_t_self0 <= 3'd6;
		end
		4'd10: begin
			builder_sync_f_t_self0 <= 2'd2;
		end
		4'd11: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
		4'd12: begin
			builder_sync_f_t_self0 <= 2'd3;
		end
		4'd13: begin
			builder_sync_f_t_self0 <= 3'd4;
		end
		4'd14: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
		default: begin
			builder_sync_f_t_self0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_303 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_304;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_self0 <= 3'd0;
	case (main_genericstandalone_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			builder_sync_f_rhs_self0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_rhs_self0 <= 3'd7;
		end
		2'd2: begin
			builder_sync_f_rhs_self0 <= 3'd4;
		end
		2'd3: begin
			builder_sync_f_rhs_self0 <= 2'd3;
		end
		3'd4: begin
			builder_sync_f_rhs_self0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_f_rhs_self0 <= 2'd2;
		end
		3'd6: begin
			builder_sync_f_rhs_self0 <= 3'd6;
		end
		3'd7: begin
			builder_sync_f_rhs_self0 <= 3'd7;
		end
		4'd8: begin
			builder_sync_f_rhs_self0 <= 3'd7;
		end
		4'd9: begin
			builder_sync_f_rhs_self0 <= 1'd1;
		end
		4'd10: begin
			builder_sync_f_rhs_self0 <= 3'd5;
		end
		4'd11: begin
			builder_sync_f_rhs_self0 <= 1'd0;
		end
		4'd12: begin
			builder_sync_f_rhs_self0 <= 2'd3;
		end
		4'd13: begin
			builder_sync_f_rhs_self0 <= 3'd4;
		end
		4'd14: begin
			builder_sync_f_rhs_self0 <= 3'd7;
		end
		default: begin
			builder_sync_f_rhs_self0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_304 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_305;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_self0 <= 5'd0;
	case (main_genericstandalone_pcs_receivepath_input_msb_first[9:4])
		1'd0: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		2'd2: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		2'd3: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		3'd4: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_rhs_self0 <= 5'd23;
		end
		3'd6: begin
			builder_sync_rhs_self0 <= 4'd8;
		end
		3'd7: begin
			builder_sync_rhs_self0 <= 3'd7;
		end
		4'd8: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		4'd9: begin
			builder_sync_rhs_self0 <= 5'd27;
		end
		4'd10: begin
			builder_sync_rhs_self0 <= 3'd4;
		end
		4'd11: begin
			builder_sync_rhs_self0 <= 5'd20;
		end
		4'd12: begin
			builder_sync_rhs_self0 <= 5'd24;
		end
		4'd13: begin
			builder_sync_rhs_self0 <= 4'd12;
		end
		4'd14: begin
			builder_sync_rhs_self0 <= 5'd28;
		end
		4'd15: begin
			builder_sync_rhs_self0 <= 5'd28;
		end
		5'd16: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		5'd17: begin
			builder_sync_rhs_self0 <= 5'd29;
		end
		5'd18: begin
			builder_sync_rhs_self0 <= 2'd2;
		end
		5'd19: begin
			builder_sync_rhs_self0 <= 5'd18;
		end
		5'd20: begin
			builder_sync_rhs_self0 <= 5'd31;
		end
		5'd21: begin
			builder_sync_rhs_self0 <= 4'd10;
		end
		5'd22: begin
			builder_sync_rhs_self0 <= 5'd26;
		end
		5'd23: begin
			builder_sync_rhs_self0 <= 4'd15;
		end
		5'd24: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		5'd25: begin
			builder_sync_rhs_self0 <= 3'd6;
		end
		5'd26: begin
			builder_sync_rhs_self0 <= 5'd22;
		end
		5'd27: begin
			builder_sync_rhs_self0 <= 5'd16;
		end
		5'd28: begin
			builder_sync_rhs_self0 <= 4'd14;
		end
		5'd29: begin
			builder_sync_rhs_self0 <= 1'd1;
		end
		5'd30: begin
			builder_sync_rhs_self0 <= 5'd30;
		end
		5'd31: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		6'd32: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		6'd33: begin
			builder_sync_rhs_self0 <= 5'd30;
		end
		6'd34: begin
			builder_sync_rhs_self0 <= 1'd1;
		end
		6'd35: begin
			builder_sync_rhs_self0 <= 5'd17;
		end
		6'd36: begin
			builder_sync_rhs_self0 <= 5'd16;
		end
		6'd37: begin
			builder_sync_rhs_self0 <= 4'd9;
		end
		6'd38: begin
			builder_sync_rhs_self0 <= 5'd25;
		end
		6'd39: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		6'd40: begin
			builder_sync_rhs_self0 <= 4'd15;
		end
		6'd41: begin
			builder_sync_rhs_self0 <= 3'd5;
		end
		6'd42: begin
			builder_sync_rhs_self0 <= 5'd21;
		end
		6'd43: begin
			builder_sync_rhs_self0 <= 5'd31;
		end
		6'd44: begin
			builder_sync_rhs_self0 <= 4'd13;
		end
		6'd45: begin
			builder_sync_rhs_self0 <= 2'd2;
		end
		6'd46: begin
			builder_sync_rhs_self0 <= 5'd29;
		end
		6'd47: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		6'd48: begin
			builder_sync_rhs_self0 <= 5'd28;
		end
		6'd49: begin
			builder_sync_rhs_self0 <= 2'd3;
		end
		6'd50: begin
			builder_sync_rhs_self0 <= 5'd19;
		end
		6'd51: begin
			builder_sync_rhs_self0 <= 5'd24;
		end
		6'd52: begin
			builder_sync_rhs_self0 <= 4'd11;
		end
		6'd53: begin
			builder_sync_rhs_self0 <= 3'd4;
		end
		6'd54: begin
			builder_sync_rhs_self0 <= 5'd27;
		end
		6'd55: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		6'd56: begin
			builder_sync_rhs_self0 <= 3'd7;
		end
		6'd57: begin
			builder_sync_rhs_self0 <= 4'd8;
		end
		6'd58: begin
			builder_sync_rhs_self0 <= 5'd23;
		end
		6'd59: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		6'd60: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		6'd61: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		6'd62: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
		default: begin
			builder_sync_rhs_self0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_305 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_306;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_self1 <= 6'd0;
	case (main_genericstandalone_pcs_transmitpath_encoder_d[4:0])
		1'd0: begin
			builder_sync_f_rhs_self1 <= 5'd24;
		end
		1'd1: begin
			builder_sync_f_rhs_self1 <= 6'd34;
		end
		2'd2: begin
			builder_sync_f_rhs_self1 <= 5'd18;
		end
		2'd3: begin
			builder_sync_f_rhs_self1 <= 6'd49;
		end
		3'd4: begin
			builder_sync_f_rhs_self1 <= 4'd10;
		end
		3'd5: begin
			builder_sync_f_rhs_self1 <= 6'd41;
		end
		3'd6: begin
			builder_sync_f_rhs_self1 <= 5'd25;
		end
		3'd7: begin
			builder_sync_f_rhs_self1 <= 3'd7;
		end
		4'd8: begin
			builder_sync_f_rhs_self1 <= 3'd6;
		end
		4'd9: begin
			builder_sync_f_rhs_self1 <= 6'd37;
		end
		4'd10: begin
			builder_sync_f_rhs_self1 <= 5'd21;
		end
		4'd11: begin
			builder_sync_f_rhs_self1 <= 6'd52;
		end
		4'd12: begin
			builder_sync_f_rhs_self1 <= 4'd13;
		end
		4'd13: begin
			builder_sync_f_rhs_self1 <= 6'd44;
		end
		4'd14: begin
			builder_sync_f_rhs_self1 <= 5'd28;
		end
		4'd15: begin
			builder_sync_f_rhs_self1 <= 6'd40;
		end
		5'd16: begin
			builder_sync_f_rhs_self1 <= 6'd36;
		end
		5'd17: begin
			builder_sync_f_rhs_self1 <= 6'd35;
		end
		5'd18: begin
			builder_sync_f_rhs_self1 <= 5'd19;
		end
		5'd19: begin
			builder_sync_f_rhs_self1 <= 6'd50;
		end
		5'd20: begin
			builder_sync_f_rhs_self1 <= 4'd11;
		end
		5'd21: begin
			builder_sync_f_rhs_self1 <= 6'd42;
		end
		5'd22: begin
			builder_sync_f_rhs_self1 <= 5'd26;
		end
		5'd23: begin
			builder_sync_f_rhs_self1 <= 3'd5;
		end
		5'd24: begin
			builder_sync_f_rhs_self1 <= 4'd12;
		end
		5'd25: begin
			builder_sync_f_rhs_self1 <= 6'd38;
		end
		5'd26: begin
			builder_sync_f_rhs_self1 <= 5'd22;
		end
		5'd27: begin
			builder_sync_f_rhs_self1 <= 4'd9;
		end
		5'd28: begin
			builder_sync_f_rhs_self1 <= 4'd14;
		end
		5'd29: begin
			builder_sync_f_rhs_self1 <= 5'd17;
		end
		5'd30: begin
			builder_sync_f_rhs_self1 <= 6'd33;
		end
		default: begin
			builder_sync_f_rhs_self1 <= 5'd20;
		end
	endcase
// synthesis translate_off
	dummy_d_306 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_307;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_self2 <= 1'd0;
	case (main_genericstandalone_pcs_transmitpath_encoder_d[4:0])
		1'd0: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		1'd1: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		2'd3: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		3'd4: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		3'd5: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		3'd6: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		3'd7: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		4'd8: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		4'd9: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		4'd10: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		4'd11: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		4'd12: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		4'd13: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		4'd14: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		4'd15: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		5'd16: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		5'd17: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd18: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd19: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd20: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd21: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd22: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd23: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		5'd24: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		5'd25: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd26: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd27: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		5'd28: begin
			builder_sync_f_rhs_self2 <= 1'd0;
		end
		5'd29: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		5'd30: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
		default: begin
			builder_sync_f_rhs_self2 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_307 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_308;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_self3 <= 1'd0;
	case (main_genericstandalone_pcs_transmitpath_encoder_d[4:0])
		1'd0: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		1'd1: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		2'd3: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		3'd4: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		3'd5: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		3'd6: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		3'd7: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		4'd8: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		4'd9: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		4'd10: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		4'd11: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		4'd12: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		4'd13: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		4'd14: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		4'd15: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		5'd16: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		5'd17: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd18: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd19: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd20: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd21: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd22: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd23: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		5'd24: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		5'd25: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd26: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd27: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		5'd28: begin
			builder_sync_f_rhs_self3 <= 1'd0;
		end
		5'd29: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		5'd30: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
		default: begin
			builder_sync_f_rhs_self3 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_308 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_309;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_self1 <= 4'd0;
	case (main_genericstandalone_pcs_transmitpath_encoder_d[7:5])
		1'd0: begin
			builder_sync_rhs_self1 <= 3'd4;
		end
		1'd1: begin
			builder_sync_rhs_self1 <= 4'd9;
		end
		2'd2: begin
			builder_sync_rhs_self1 <= 3'd5;
		end
		2'd3: begin
			builder_sync_rhs_self1 <= 2'd3;
		end
		3'd4: begin
			builder_sync_rhs_self1 <= 2'd2;
		end
		3'd5: begin
			builder_sync_rhs_self1 <= 4'd10;
		end
		3'd6: begin
			builder_sync_rhs_self1 <= 3'd6;
		end
		default: begin
			builder_sync_rhs_self1 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_309 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_310;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_self2 <= 1'd0;
	case (main_genericstandalone_pcs_transmitpath_encoder_d[7:5])
		1'd0: begin
			builder_sync_rhs_self2 <= 1'd1;
		end
		1'd1: begin
			builder_sync_rhs_self2 <= 1'd0;
		end
		2'd2: begin
			builder_sync_rhs_self2 <= 1'd0;
		end
		2'd3: begin
			builder_sync_rhs_self2 <= 1'd0;
		end
		3'd4: begin
			builder_sync_rhs_self2 <= 1'd1;
		end
		3'd5: begin
			builder_sync_rhs_self2 <= 1'd0;
		end
		3'd6: begin
			builder_sync_rhs_self2 <= 1'd0;
		end
		default: begin
			builder_sync_rhs_self2 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_310 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_311;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_self4 <= 1'd0;
	case (main_genericstandalone_pcs_transmitpath_encoder_d[7:5])
		1'd0: begin
			builder_sync_f_rhs_self4 <= 1'd1;
		end
		1'd1: begin
			builder_sync_f_rhs_self4 <= 1'd0;
		end
		2'd2: begin
			builder_sync_f_rhs_self4 <= 1'd0;
		end
		2'd3: begin
			builder_sync_f_rhs_self4 <= 1'd1;
		end
		3'd4: begin
			builder_sync_f_rhs_self4 <= 1'd1;
		end
		3'd5: begin
			builder_sync_f_rhs_self4 <= 1'd0;
		end
		3'd6: begin
			builder_sync_f_rhs_self4 <= 1'd0;
		end
		default: begin
			builder_sync_f_rhs_self4 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_311 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_312;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_self3 <= 61'd0;
	case (main_genericstandalone_rtio_core_sed_lane_dist_current_lane)
		1'd0: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps0;
		end
		1'd1: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps1;
		end
		2'd2: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps2;
		end
		2'd3: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps3;
		end
		3'd4: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps4;
		end
		3'd5: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps5;
		end
		3'd6: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps6;
		end
		3'd7: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps7;
		end
		4'd8: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps8;
		end
		4'd9: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps9;
		end
		4'd10: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps10;
		end
		4'd11: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps11;
		end
		4'd12: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps12;
		end
		4'd13: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps13;
		end
		4'd14: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps14;
		end
		default: begin
			builder_sync_rhs_self3 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps15;
		end
	endcase
// synthesis translate_off
	dummy_d_312 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_313;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_self4 <= 61'd0;
	case (main_genericstandalone_rtio_core_sed_lane_dist_current_lane_plus_one)
		1'd0: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps0;
		end
		1'd1: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps1;
		end
		2'd2: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps2;
		end
		2'd3: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps3;
		end
		3'd4: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps4;
		end
		3'd5: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps5;
		end
		3'd6: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps6;
		end
		3'd7: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps7;
		end
		4'd8: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps8;
		end
		4'd9: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps9;
		end
		4'd10: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps10;
		end
		4'd11: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps11;
		end
		4'd12: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps12;
		end
		4'd13: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps13;
		end
		4'd14: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps14;
		end
		default: begin
			builder_sync_rhs_self4 <= main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps15;
		end
	endcase
// synthesis translate_off
	dummy_d_313 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_314;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self0 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r0)
		1'd0: begin
			builder_sync_basiclowerer_self0 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self0 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self0 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self0 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self0 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self0 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self0 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self0 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self0 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self0 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self0 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self0 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self0 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self0 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self0 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self0 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self0 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self0 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self0 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self0 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self0 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self0 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self0 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self0 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self0 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self0 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self0 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self0 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self0 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self0 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self0 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self0 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self0 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self0 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self0 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self0 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self0 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self0 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_314 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_315;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self1 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r1)
		1'd0: begin
			builder_sync_basiclowerer_self1 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self1 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self1 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self1 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self1 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self1 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self1 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self1 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self1 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self1 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self1 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self1 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self1 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self1 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self1 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self1 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self1 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self1 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self1 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self1 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self1 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self1 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self1 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self1 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self1 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self1 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self1 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self1 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self1 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self1 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self1 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self1 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self1 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self1 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self1 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self1 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self1 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self1 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_315 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_316;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self2 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r2)
		1'd0: begin
			builder_sync_basiclowerer_self2 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self2 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self2 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self2 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self2 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self2 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self2 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self2 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self2 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self2 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self2 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self2 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self2 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self2 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self2 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self2 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self2 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self2 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self2 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self2 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self2 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self2 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self2 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self2 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self2 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self2 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self2 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self2 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self2 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self2 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self2 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self2 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self2 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self2 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self2 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self2 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self2 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self2 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_316 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_317;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self3 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r3)
		1'd0: begin
			builder_sync_basiclowerer_self3 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self3 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self3 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self3 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self3 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self3 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self3 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self3 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self3 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self3 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self3 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self3 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self3 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self3 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self3 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self3 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self3 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self3 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self3 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self3 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self3 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self3 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self3 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self3 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self3 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self3 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self3 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self3 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self3 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self3 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self3 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self3 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self3 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self3 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self3 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self3 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self3 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self3 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_317 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_318;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self4 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r4)
		1'd0: begin
			builder_sync_basiclowerer_self4 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self4 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self4 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self4 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self4 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self4 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self4 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self4 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self4 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self4 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self4 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self4 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self4 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self4 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self4 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self4 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self4 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self4 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self4 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self4 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self4 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self4 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self4 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self4 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self4 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self4 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self4 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self4 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self4 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self4 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self4 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self4 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self4 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self4 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self4 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self4 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self4 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self4 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_318 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_319;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self5 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r5)
		1'd0: begin
			builder_sync_basiclowerer_self5 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self5 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self5 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self5 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self5 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self5 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self5 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self5 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self5 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self5 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self5 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self5 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self5 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self5 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self5 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self5 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self5 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self5 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self5 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self5 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self5 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self5 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self5 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self5 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self5 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self5 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self5 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self5 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self5 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self5 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self5 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self5 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self5 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self5 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self5 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self5 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self5 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self5 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_319 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_320;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self6 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r6)
		1'd0: begin
			builder_sync_basiclowerer_self6 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self6 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self6 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self6 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self6 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self6 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self6 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self6 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self6 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self6 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self6 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self6 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self6 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self6 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self6 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self6 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self6 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self6 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self6 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self6 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self6 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self6 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self6 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self6 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self6 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self6 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self6 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self6 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self6 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self6 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self6 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self6 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self6 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self6 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self6 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self6 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self6 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self6 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_320 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_321;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self7 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r7)
		1'd0: begin
			builder_sync_basiclowerer_self7 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self7 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self7 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self7 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self7 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self7 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self7 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self7 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self7 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self7 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self7 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self7 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self7 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self7 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self7 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self7 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self7 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self7 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self7 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self7 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self7 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self7 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self7 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self7 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self7 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self7 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self7 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self7 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self7 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self7 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self7 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self7 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self7 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self7 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self7 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self7 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self7 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self7 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_321 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_322;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self8 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r8)
		1'd0: begin
			builder_sync_basiclowerer_self8 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self8 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self8 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self8 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self8 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self8 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self8 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self8 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self8 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self8 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self8 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self8 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self8 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self8 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self8 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self8 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self8 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self8 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self8 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self8 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self8 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self8 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self8 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self8 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self8 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self8 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self8 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self8 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self8 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self8 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self8 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self8 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self8 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self8 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self8 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self8 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self8 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self8 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_322 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_323;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self9 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r9)
		1'd0: begin
			builder_sync_basiclowerer_self9 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self9 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self9 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self9 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self9 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self9 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self9 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self9 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self9 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self9 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self9 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self9 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self9 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self9 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self9 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self9 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self9 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self9 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self9 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self9 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self9 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self9 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self9 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self9 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self9 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self9 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self9 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self9 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self9 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self9 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self9 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self9 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self9 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self9 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self9 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self9 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self9 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self9 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_323 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_324;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self10 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r10)
		1'd0: begin
			builder_sync_basiclowerer_self10 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self10 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self10 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self10 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self10 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self10 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self10 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self10 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self10 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self10 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self10 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self10 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self10 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self10 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self10 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self10 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self10 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self10 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self10 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self10 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self10 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self10 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self10 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self10 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self10 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self10 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self10 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self10 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self10 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self10 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self10 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self10 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self10 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self10 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self10 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self10 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self10 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self10 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_324 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_325;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self11 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r11)
		1'd0: begin
			builder_sync_basiclowerer_self11 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self11 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self11 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self11 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self11 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self11 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self11 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self11 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self11 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self11 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self11 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self11 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self11 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self11 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self11 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self11 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self11 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self11 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self11 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self11 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self11 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self11 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self11 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self11 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self11 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self11 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self11 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self11 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self11 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self11 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self11 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self11 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self11 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self11 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self11 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self11 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self11 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self11 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_325 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_326;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self12 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r12)
		1'd0: begin
			builder_sync_basiclowerer_self12 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self12 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self12 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self12 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self12 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self12 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self12 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self12 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self12 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self12 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self12 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self12 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self12 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self12 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self12 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self12 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self12 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self12 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self12 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self12 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self12 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self12 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self12 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self12 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self12 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self12 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self12 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self12 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self12 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self12 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self12 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self12 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self12 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self12 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self12 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self12 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self12 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self12 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_326 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_327;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self13 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r13)
		1'd0: begin
			builder_sync_basiclowerer_self13 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self13 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self13 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self13 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self13 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self13 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self13 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self13 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self13 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self13 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self13 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self13 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self13 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self13 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self13 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self13 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self13 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self13 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self13 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self13 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self13 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self13 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self13 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self13 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self13 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self13 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self13 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self13 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self13 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self13 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self13 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self13 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self13 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self13 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self13 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self13 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self13 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self13 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_327 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_328;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self14 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r14)
		1'd0: begin
			builder_sync_basiclowerer_self14 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self14 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self14 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self14 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self14 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self14 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self14 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self14 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self14 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self14 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self14 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self14 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self14 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self14 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self14 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self14 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self14 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self14 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self14 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self14 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self14 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self14 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self14 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self14 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self14 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self14 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self14 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self14 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self14 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self14 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self14 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self14 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self14 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self14 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self14 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self14 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self14 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self14 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_328 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_329;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_self15 <= 1'd0;
	case (main_genericstandalone_rtio_core_sed_channel_r15)
		1'd0: begin
			builder_sync_basiclowerer_self15 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_self15 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_self15 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_self15 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_self15 <= main_output_8x0_busy0;
		end
		3'd5: begin
			builder_sync_basiclowerer_self15 <= main_output_8x1_busy0;
		end
		3'd6: begin
			builder_sync_basiclowerer_self15 <= main_output_8x2_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_self15 <= main_output_8x3_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_self15 <= main_output_8x4_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_self15 <= main_output_8x5_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_self15 <= main_output_8x6_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_self15 <= main_output_8x7_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_self15 <= main_output_8x8_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_self15 <= main_output_8x9_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_self15 <= main_output_8x10_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_self15 <= main_output_8x11_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_self15 <= main_spimaster0_ointerface0_busy0;
		end
		5'd17: begin
			builder_sync_basiclowerer_self15 <= main_output_8x0_busy1;
		end
		5'd18: begin
			builder_sync_basiclowerer_self15 <= main_output_8x12_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_self15 <= main_output_8x13_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_self15 <= main_output_8x14_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_self15 <= main_output_8x15_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_self15 <= main_spimaster1_ointerface1_busy0;
		end
		5'd23: begin
			builder_sync_basiclowerer_self15 <= main_output_8x1_busy1;
		end
		5'd24: begin
			builder_sync_basiclowerer_self15 <= main_output_8x16_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_self15 <= main_output_8x17_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_self15 <= main_output_8x18_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_self15 <= main_output_8x19_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_self15 <= main_spimaster0_ointerface0_busy1;
		end
		5'd29: begin
			builder_sync_basiclowerer_self15 <= main_spimaster1_ointerface1_busy1;
		end
		5'd30: begin
			builder_sync_basiclowerer_self15 <= main_output_8x20_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_self15 <= main_spimaster2_ointerface2_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_self15 <= main_ldac_phy_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_self15 <= main_clr_phy_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_self15 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_self15 <= main_output1_busy;
		end
		6'd36: begin
			builder_sync_basiclowerer_self15 <= main_output2_busy;
		end
		default: begin
			builder_sync_basiclowerer_self15 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_329 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_330;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self1 <= 32'd0;
	case (main_genericstandalone_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record0_fifo_out_data;
		end
		1'd1: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record1_fifo_out_data;
		end
		2'd2: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record2_fifo_out_data;
		end
		2'd3: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record3_fifo_out_data;
		end
		3'd4: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record4_fifo_out_data;
		end
		5'd17: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record5_fifo_out_data;
		end
		5'd23: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record6_fifo_out_data;
		end
		5'd29: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record7_fifo_out_data;
		end
		5'd30: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		5'd31: begin
			builder_sync_t_rhs_self1 <= main_genericstandalone_rtio_core_inputcollector_record8_fifo_out_data;
		end
		6'd32: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		6'd33: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		6'd34: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		6'd35: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		6'd36: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self1 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_330 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_331;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self2 <= 65'd0;
	case (main_genericstandalone_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_sync_t_rhs_self2 <= (main_genericstandalone_rtio_core_inputcollector_record0_fifo_out_timestamp <<< 1'd0);
		end
		1'd1: begin
			builder_sync_t_rhs_self2 <= (main_genericstandalone_rtio_core_inputcollector_record1_fifo_out_timestamp <<< 1'd0);
		end
		2'd2: begin
			builder_sync_t_rhs_self2 <= (main_genericstandalone_rtio_core_inputcollector_record2_fifo_out_timestamp <<< 1'd0);
		end
		2'd3: begin
			builder_sync_t_rhs_self2 <= (main_genericstandalone_rtio_core_inputcollector_record3_fifo_out_timestamp <<< 1'd0);
		end
		3'd4: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		5'd31: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		6'd32: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		6'd33: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		6'd34: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		6'd35: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		6'd36: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self2 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_331 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_332;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self1 <= 8'd0;
	case (main_inout_8x0_inout_8x0_ointerface0_fine_ts)
		1'd0: begin
			builder_sync_f_t_self1 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self1 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self1 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self1 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self1 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self1 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self1 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self1 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_332 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_333;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self2 <= 7'd0;
	case (main_inout_8x0_inout_8x0_ointerface0_fine_ts)
		1'd0: begin
			builder_sync_f_t_self2 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self2 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self2 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self2 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self2 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self2 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self2 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self2 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_333 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_334;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self3 <= 8'd0;
	case (main_inout_8x1_inout_8x1_ointerface1_fine_ts)
		1'd0: begin
			builder_sync_f_t_self3 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self3 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self3 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self3 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self3 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self3 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self3 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self3 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_334 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_335;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self4 <= 7'd0;
	case (main_inout_8x1_inout_8x1_ointerface1_fine_ts)
		1'd0: begin
			builder_sync_f_t_self4 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self4 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self4 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self4 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self4 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self4 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self4 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self4 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_335 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_336;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self5 <= 8'd0;
	case (main_inout_8x2_inout_8x2_ointerface2_fine_ts)
		1'd0: begin
			builder_sync_f_t_self5 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self5 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self5 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self5 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self5 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self5 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self5 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self5 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_336 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_337;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self6 <= 7'd0;
	case (main_inout_8x2_inout_8x2_ointerface2_fine_ts)
		1'd0: begin
			builder_sync_f_t_self6 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self6 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self6 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self6 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self6 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self6 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self6 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self6 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_337 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_338;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self7 <= 8'd0;
	case (main_inout_8x3_inout_8x3_ointerface3_fine_ts)
		1'd0: begin
			builder_sync_f_t_self7 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self7 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self7 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self7 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self7 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self7 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self7 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self7 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_338 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_339;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self8 <= 7'd0;
	case (main_inout_8x3_inout_8x3_ointerface3_fine_ts)
		1'd0: begin
			builder_sync_f_t_self8 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self8 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self8 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self8 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self8 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self8 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self8 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self8 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_339 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_340;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self9 <= 8'd0;
	case (main_output_8x0_fine_ts0)
		1'd0: begin
			builder_sync_f_t_self9 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self9 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self9 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self9 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self9 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self9 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self9 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self9 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_340 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_341;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self10 <= 7'd0;
	case (main_output_8x0_fine_ts0)
		1'd0: begin
			builder_sync_f_t_self10 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self10 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self10 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self10 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self10 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self10 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self10 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self10 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_341 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_342;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self11 <= 8'd0;
	case (main_output_8x1_fine_ts0)
		1'd0: begin
			builder_sync_f_t_self11 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self11 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self11 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self11 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self11 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self11 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self11 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self11 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_342 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_343;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self12 <= 7'd0;
	case (main_output_8x1_fine_ts0)
		1'd0: begin
			builder_sync_f_t_self12 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self12 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self12 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self12 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self12 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self12 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self12 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self12 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_343 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_344;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self13 <= 8'd0;
	case (main_output_8x2_fine_ts)
		1'd0: begin
			builder_sync_f_t_self13 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self13 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self13 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self13 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self13 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self13 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self13 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self13 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_344 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_345;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self14 <= 7'd0;
	case (main_output_8x2_fine_ts)
		1'd0: begin
			builder_sync_f_t_self14 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self14 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self14 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self14 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self14 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self14 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self14 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self14 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_345 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_346;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self15 <= 8'd0;
	case (main_output_8x3_fine_ts)
		1'd0: begin
			builder_sync_f_t_self15 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self15 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self15 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self15 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self15 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self15 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self15 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self15 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_346 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_347;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self16 <= 7'd0;
	case (main_output_8x3_fine_ts)
		1'd0: begin
			builder_sync_f_t_self16 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self16 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self16 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self16 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self16 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self16 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self16 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self16 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_347 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_348;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self17 <= 8'd0;
	case (main_output_8x4_fine_ts)
		1'd0: begin
			builder_sync_f_t_self17 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self17 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self17 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self17 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self17 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self17 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self17 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self17 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_348 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_349;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self18 <= 7'd0;
	case (main_output_8x4_fine_ts)
		1'd0: begin
			builder_sync_f_t_self18 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self18 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self18 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self18 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self18 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self18 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self18 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self18 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_349 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_350;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self19 <= 8'd0;
	case (main_output_8x5_fine_ts)
		1'd0: begin
			builder_sync_f_t_self19 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self19 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self19 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self19 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self19 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self19 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self19 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self19 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_350 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_351;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self20 <= 7'd0;
	case (main_output_8x5_fine_ts)
		1'd0: begin
			builder_sync_f_t_self20 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self20 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self20 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self20 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self20 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self20 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self20 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self20 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_351 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_352;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self21 <= 8'd0;
	case (main_output_8x6_fine_ts)
		1'd0: begin
			builder_sync_f_t_self21 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self21 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self21 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self21 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self21 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self21 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self21 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self21 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_352 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_353;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self22 <= 7'd0;
	case (main_output_8x6_fine_ts)
		1'd0: begin
			builder_sync_f_t_self22 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self22 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self22 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self22 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self22 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self22 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self22 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self22 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_353 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_354;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self23 <= 8'd0;
	case (main_output_8x7_fine_ts)
		1'd0: begin
			builder_sync_f_t_self23 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self23 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self23 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self23 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self23 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self23 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self23 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self23 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_354 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_355;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self24 <= 7'd0;
	case (main_output_8x7_fine_ts)
		1'd0: begin
			builder_sync_f_t_self24 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self24 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self24 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self24 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self24 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self24 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self24 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self24 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_355 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_356;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self25 <= 8'd0;
	case (main_output_8x8_fine_ts)
		1'd0: begin
			builder_sync_f_t_self25 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self25 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self25 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self25 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self25 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self25 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self25 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self25 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_356 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_357;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self26 <= 7'd0;
	case (main_output_8x8_fine_ts)
		1'd0: begin
			builder_sync_f_t_self26 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self26 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self26 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self26 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self26 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self26 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self26 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self26 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_357 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_358;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self27 <= 8'd0;
	case (main_output_8x9_fine_ts)
		1'd0: begin
			builder_sync_f_t_self27 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self27 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self27 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self27 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self27 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self27 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self27 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self27 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_358 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_359;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self28 <= 7'd0;
	case (main_output_8x9_fine_ts)
		1'd0: begin
			builder_sync_f_t_self28 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self28 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self28 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self28 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self28 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self28 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self28 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self28 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_359 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_360;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self29 <= 8'd0;
	case (main_output_8x10_fine_ts)
		1'd0: begin
			builder_sync_f_t_self29 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self29 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self29 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self29 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self29 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self29 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self29 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self29 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_360 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_361;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self30 <= 7'd0;
	case (main_output_8x10_fine_ts)
		1'd0: begin
			builder_sync_f_t_self30 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self30 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self30 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self30 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self30 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self30 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self30 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self30 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_361 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_362;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self31 <= 8'd0;
	case (main_output_8x11_fine_ts)
		1'd0: begin
			builder_sync_f_t_self31 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self31 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self31 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self31 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self31 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self31 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self31 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self31 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_362 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_363;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self32 <= 7'd0;
	case (main_output_8x11_fine_ts)
		1'd0: begin
			builder_sync_f_t_self32 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self32 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self32 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self32 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self32 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self32 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self32 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self32 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_363 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_364;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self33 <= 8'd0;
	case (main_output_8x0_fine_ts1)
		1'd0: begin
			builder_sync_f_t_self33 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self33 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self33 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self33 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self33 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self33 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self33 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self33 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_364 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_365;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self34 <= 7'd0;
	case (main_output_8x0_fine_ts1)
		1'd0: begin
			builder_sync_f_t_self34 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self34 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self34 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self34 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self34 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self34 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self34 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self34 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_365 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_366;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self35 <= 8'd0;
	case (main_output_8x12_fine_ts)
		1'd0: begin
			builder_sync_f_t_self35 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self35 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self35 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self35 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self35 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self35 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self35 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self35 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_366 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_367;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self36 <= 7'd0;
	case (main_output_8x12_fine_ts)
		1'd0: begin
			builder_sync_f_t_self36 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self36 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self36 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self36 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self36 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self36 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self36 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self36 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_367 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_368;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self37 <= 8'd0;
	case (main_output_8x13_fine_ts)
		1'd0: begin
			builder_sync_f_t_self37 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self37 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self37 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self37 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self37 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self37 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self37 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self37 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_368 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_369;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self38 <= 7'd0;
	case (main_output_8x13_fine_ts)
		1'd0: begin
			builder_sync_f_t_self38 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self38 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self38 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self38 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self38 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self38 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self38 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self38 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_369 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_370;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self39 <= 8'd0;
	case (main_output_8x14_fine_ts)
		1'd0: begin
			builder_sync_f_t_self39 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self39 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self39 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self39 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self39 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self39 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self39 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self39 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_370 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_371;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self40 <= 7'd0;
	case (main_output_8x14_fine_ts)
		1'd0: begin
			builder_sync_f_t_self40 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self40 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self40 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self40 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self40 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self40 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self40 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self40 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_371 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_372;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self41 <= 8'd0;
	case (main_output_8x15_fine_ts)
		1'd0: begin
			builder_sync_f_t_self41 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self41 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self41 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self41 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self41 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self41 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self41 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self41 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_372 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_373;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self42 <= 7'd0;
	case (main_output_8x15_fine_ts)
		1'd0: begin
			builder_sync_f_t_self42 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self42 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self42 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self42 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self42 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self42 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self42 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self42 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_373 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_374;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self43 <= 8'd0;
	case (main_output_8x1_fine_ts1)
		1'd0: begin
			builder_sync_f_t_self43 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self43 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self43 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self43 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self43 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self43 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self43 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self43 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_374 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_375;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self44 <= 7'd0;
	case (main_output_8x1_fine_ts1)
		1'd0: begin
			builder_sync_f_t_self44 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self44 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self44 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self44 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self44 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self44 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self44 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self44 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_375 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_376;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self45 <= 8'd0;
	case (main_output_8x16_fine_ts)
		1'd0: begin
			builder_sync_f_t_self45 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self45 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self45 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self45 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self45 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self45 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self45 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self45 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_376 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_377;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self46 <= 7'd0;
	case (main_output_8x16_fine_ts)
		1'd0: begin
			builder_sync_f_t_self46 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self46 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self46 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self46 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self46 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self46 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self46 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self46 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_377 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_378;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self47 <= 8'd0;
	case (main_output_8x17_fine_ts)
		1'd0: begin
			builder_sync_f_t_self47 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self47 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self47 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self47 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self47 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self47 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self47 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self47 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_378 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_379;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self48 <= 7'd0;
	case (main_output_8x17_fine_ts)
		1'd0: begin
			builder_sync_f_t_self48 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self48 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self48 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self48 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self48 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self48 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self48 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self48 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_379 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_380;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self49 <= 8'd0;
	case (main_output_8x18_fine_ts)
		1'd0: begin
			builder_sync_f_t_self49 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self49 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self49 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self49 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self49 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self49 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self49 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self49 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_380 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_381;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self50 <= 7'd0;
	case (main_output_8x18_fine_ts)
		1'd0: begin
			builder_sync_f_t_self50 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self50 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self50 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self50 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self50 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self50 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self50 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self50 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_381 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_382;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self51 <= 8'd0;
	case (main_output_8x19_fine_ts)
		1'd0: begin
			builder_sync_f_t_self51 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self51 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self51 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self51 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self51 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self51 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self51 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self51 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_382 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_383;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self52 <= 7'd0;
	case (main_output_8x19_fine_ts)
		1'd0: begin
			builder_sync_f_t_self52 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self52 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self52 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self52 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self52 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self52 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self52 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self52 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_383 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_384;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self53 <= 8'd0;
	case (main_output_8x20_fine_ts)
		1'd0: begin
			builder_sync_f_t_self53 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self53 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self53 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self53 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self53 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self53 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self53 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self53 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_384 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_385;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self54 <= 7'd0;
	case (main_output_8x20_fine_ts)
		1'd0: begin
			builder_sync_f_t_self54 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self54 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self54 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self54 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self54 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self54 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self54 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self54 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_385 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_386;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self55 <= 8'd0;
	case (main_ldac_phy_fine_ts)
		1'd0: begin
			builder_sync_f_t_self55 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self55 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self55 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self55 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self55 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self55 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self55 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self55 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_386 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_387;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self56 <= 7'd0;
	case (main_ldac_phy_fine_ts)
		1'd0: begin
			builder_sync_f_t_self56 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self56 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self56 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self56 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self56 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self56 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self56 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self56 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_387 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_388;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self57 <= 8'd0;
	case (main_clr_phy_fine_ts)
		1'd0: begin
			builder_sync_f_t_self57 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_self57 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_self57 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_self57 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_self57 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_self57 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_self57 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_self57 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_388 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_389;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_self58 <= 7'd0;
	case (main_clr_phy_fine_ts)
		1'd0: begin
			builder_sync_f_t_self58 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_self58 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_self58 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_self58 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_self58 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_self58 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_self58 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_self58 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_389 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_390;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_self5 <= 32'd0;
	case (main_genericstandalone_mailbox_i1_adr[1:0])
		1'd0: begin
			builder_sync_rhs_self5 <= main_genericstandalone_mailbox0;
		end
		1'd1: begin
			builder_sync_rhs_self5 <= main_genericstandalone_mailbox1;
		end
		default: begin
			builder_sync_rhs_self5 <= main_genericstandalone_mailbox2;
		end
	endcase
// synthesis translate_off
	dummy_d_390 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_391;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_self6 <= 32'd0;
	case (main_genericstandalone_mailbox_i2_adr[1:0])
		1'd0: begin
			builder_sync_rhs_self6 <= main_genericstandalone_mailbox0;
		end
		1'd1: begin
			builder_sync_rhs_self6 <= main_genericstandalone_mailbox1;
		end
		default: begin
			builder_sync_rhs_self6 <= main_genericstandalone_mailbox2;
		end
	endcase
// synthesis translate_off
	dummy_d_391 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_392;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self4 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self4 <= main_genericstandalone_mon_bussynchronizer0_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self4 <= main_genericstandalone_mon_bussynchronizer1_o;
		end
		2'd2: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self4 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_392 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_393;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self5 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self5 <= main_genericstandalone_mon_bussynchronizer2_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self5 <= main_genericstandalone_mon_bussynchronizer3_o;
		end
		2'd2: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self5 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_393 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_394;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self6 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self6 <= main_genericstandalone_mon_bussynchronizer4_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self6 <= main_genericstandalone_mon_bussynchronizer5_o;
		end
		2'd2: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self6 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_394 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_395;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self7 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self7 <= main_genericstandalone_mon_bussynchronizer6_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self7 <= main_genericstandalone_mon_bussynchronizer7_o;
		end
		2'd2: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self7 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_395 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_396;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self8 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self8 <= main_genericstandalone_mon_bussynchronizer8_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self8 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_396 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_397;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self9 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self9 <= main_genericstandalone_mon_bussynchronizer9_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self9 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_397 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_398;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self10 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self10 <= main_genericstandalone_mon_bussynchronizer10_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self10 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_398 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_399;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self11 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self11 <= main_genericstandalone_mon_bussynchronizer11_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self11 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_399 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_400;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self12 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self12 <= main_genericstandalone_mon_bussynchronizer12_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self12 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_400 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_401;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self13 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self13 <= main_genericstandalone_mon_bussynchronizer13_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self13 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_401 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_402;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self14 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self14 <= main_genericstandalone_mon_bussynchronizer14_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self14 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_402 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_403;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self15 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self15 <= main_genericstandalone_mon_bussynchronizer15_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self15 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_403 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_404;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self16 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self16 <= main_genericstandalone_mon_bussynchronizer16_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self16 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_404 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_405;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self17 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self17 <= main_genericstandalone_mon_bussynchronizer17_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self17 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_405 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_406;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self18 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self18 <= main_genericstandalone_mon_bussynchronizer18_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self18 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_406 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_407;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self19 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self19 <= main_genericstandalone_mon_bussynchronizer19_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self19 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_407 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_408;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self20 <= 32'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self20 <= main_genericstandalone_mon_bussynchronizer20_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self20 <= main_genericstandalone_mon_bussynchronizer21_o;
		end
		2'd2: begin
			builder_sync_t_rhs_self20 <= main_genericstandalone_mon_bussynchronizer22_o;
		end
		2'd3: begin
			builder_sync_t_rhs_self20 <= main_genericstandalone_mon_bussynchronizer23_o;
		end
		3'd4: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self20 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_408 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_409;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self21 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self21 <= main_genericstandalone_mon_bussynchronizer24_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self21 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_409 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_410;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self22 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self22 <= main_genericstandalone_mon_bussynchronizer25_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self22 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_410 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_411;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self23 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self23 <= main_genericstandalone_mon_bussynchronizer26_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self23 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_411 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_412;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self24 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self24 <= main_genericstandalone_mon_bussynchronizer27_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self24 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_412 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_413;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self25 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self25 <= main_genericstandalone_mon_bussynchronizer28_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self25 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_413 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_414;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self26 <= 32'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self26 <= main_genericstandalone_mon_bussynchronizer29_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self26 <= main_genericstandalone_mon_bussynchronizer30_o;
		end
		2'd2: begin
			builder_sync_t_rhs_self26 <= main_genericstandalone_mon_bussynchronizer31_o;
		end
		2'd3: begin
			builder_sync_t_rhs_self26 <= main_genericstandalone_mon_bussynchronizer32_o;
		end
		3'd4: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self26 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_414 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_415;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self27 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self27 <= main_genericstandalone_mon_bussynchronizer33_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self27 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_415 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_416;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self28 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self28 <= main_genericstandalone_mon_bussynchronizer34_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self28 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_416 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_417;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self29 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self29 <= main_genericstandalone_mon_bussynchronizer35_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self29 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_417 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_418;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self30 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self30 <= main_genericstandalone_mon_bussynchronizer36_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self30 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_418 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_419;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self31 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self31 <= main_genericstandalone_mon_bussynchronizer37_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self31 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_419 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_420;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self32 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self32 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_420 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_421;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self33 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self33 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_421 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_422;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self34 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self34 <= main_genericstandalone_mon_bussynchronizer38_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self34 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_422 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_423;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self35 <= 16'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer39_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer40_o;
		end
		2'd2: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer41_o;
		end
		2'd3: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer42_o;
		end
		3'd4: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer43_o;
		end
		3'd5: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer44_o;
		end
		3'd6: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer45_o;
		end
		3'd7: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer46_o;
		end
		4'd8: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer47_o;
		end
		4'd9: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer48_o;
		end
		4'd10: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer49_o;
		end
		4'd11: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer50_o;
		end
		4'd12: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer51_o;
		end
		4'd13: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer52_o;
		end
		4'd14: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer53_o;
		end
		4'd15: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer54_o;
		end
		5'd16: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer55_o;
		end
		5'd17: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer56_o;
		end
		5'd18: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer57_o;
		end
		5'd19: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer58_o;
		end
		5'd20: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer59_o;
		end
		5'd21: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer60_o;
		end
		5'd22: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer61_o;
		end
		5'd23: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer62_o;
		end
		5'd24: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer63_o;
		end
		5'd25: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer64_o;
		end
		5'd26: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer65_o;
		end
		5'd27: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer66_o;
		end
		5'd28: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer67_o;
		end
		5'd29: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer68_o;
		end
		5'd30: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer69_o;
		end
		default: begin
			builder_sync_t_rhs_self35 <= main_genericstandalone_mon_bussynchronizer70_o;
		end
	endcase
// synthesis translate_off
	dummy_d_423 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_424;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self36 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self36 <= main_genericstandalone_mon_bussynchronizer71_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self36 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_424 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_425;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self37 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self37 <= main_genericstandalone_mon_bussynchronizer72_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self37 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_425 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_426;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self38 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self38 <= main_genericstandalone_mon_bussynchronizer73_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self38 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_426 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_427;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self39 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self39 <= main_genericstandalone_mon_bussynchronizer74_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self39 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_427 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_428;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self40 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self40 <= main_genericstandalone_mon_bussynchronizer75_o;
		end
		1'd1: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self40 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_428 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_429;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self41 <= 1'd0;
	case (main_genericstandalone_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_self41 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_429 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_430;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_self3 <= 32'd0;
	case (main_genericstandalone_mon_chan_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self4;
		end
		1'd1: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self5;
		end
		2'd2: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self6;
		end
		2'd3: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self7;
		end
		3'd4: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self8;
		end
		3'd5: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self9;
		end
		3'd6: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self10;
		end
		3'd7: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self11;
		end
		4'd8: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self12;
		end
		4'd9: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self13;
		end
		4'd10: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self14;
		end
		4'd11: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self15;
		end
		4'd12: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self16;
		end
		4'd13: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self17;
		end
		4'd14: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self18;
		end
		4'd15: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self19;
		end
		5'd16: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self20;
		end
		5'd17: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self21;
		end
		5'd18: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self22;
		end
		5'd19: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self23;
		end
		5'd20: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self24;
		end
		5'd21: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self25;
		end
		5'd22: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self26;
		end
		5'd23: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self27;
		end
		5'd24: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self28;
		end
		5'd25: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self29;
		end
		5'd26: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self30;
		end
		5'd27: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self31;
		end
		5'd28: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self32;
		end
		5'd29: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self33;
		end
		5'd30: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self34;
		end
		5'd31: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self35;
		end
		6'd32: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self36;
		end
		6'd33: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self37;
		end
		6'd34: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self38;
		end
		6'd35: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self39;
		end
		6'd36: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self40;
		end
		default: begin
			builder_sync_t_rhs_self3 <= builder_sync_t_rhs_self41;
		end
	endcase
// synthesis translate_off
	dummy_d_430 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx = builder_xilinxmultiregimpl01;
assign main_genericstandalone_genericstandalone_crg_i_switch = builder_xilinxmultiregimpl11;
assign builder_xilinxasyncresetsynchronizerimpl0_async_reset = (~main_genericstandalone_genericstandalone_crg_pll_locked);
assign main_genericstandalone_genericstandalone_crg_status = builder_xilinxmultiregimpl21;
assign main_genericstandalone_genericstandalone_icap_toggle_o = builder_xilinxmultiregimpl31;
assign main_genericstandalone_pcs_lp_abi_ping_toggle_o = builder_xilinxmultiregimpl41;
assign main_genericstandalone_pcs_lp_abi_pong_toggle_o = builder_xilinxmultiregimpl51;
assign main_genericstandalone_pcs_lp_abi_obuffer = builder_xilinxmultiregimpl61;
assign main_genericstandalone_pcs_seen_valid_ci_toggle_o = builder_xilinxmultiregimpl71;
assign main_genericstandalone_pcs_rx_config_reg_abi_toggle_o = builder_xilinxmultiregimpl81;
assign main_genericstandalone_pcs_rx_config_reg_ack_toggle_o = builder_xilinxmultiregimpl91;
assign builder_xilinxasyncresetsynchronizerimpl1_async_reset = (~main_genericstandalone_tx_mmcm_locked);
assign builder_xilinxasyncresetsynchronizerimpl2_async_reset = (~main_genericstandalone_rx_mmcm_locked);
assign main_genericstandalone_tx_init_qpll_lock1 = builder_xilinxmultiregimpl101;
assign main_genericstandalone_rx_init_rx_pma_reset_done1 = builder_xilinxmultiregimpl111;
assign main_genericstandalone_toggle_o = builder_xilinxmultiregimpl121;
assign main_genericstandalone_ps_preamble_error_toggle_o = builder_xilinxmultiregimpl131;
assign main_genericstandalone_ps_crc_error_toggle_o = builder_xilinxmultiregimpl141;
assign main_genericstandalone_tx_cdc_produce_rdomain = builder_xilinxmultiregimpl151;
assign main_genericstandalone_tx_cdc_consume_wdomain = builder_xilinxmultiregimpl161;
assign main_genericstandalone_rx_cdc_produce_rdomain = builder_xilinxmultiregimpl171;
assign main_genericstandalone_rx_cdc_consume_wdomain = builder_xilinxmultiregimpl181;
assign main_genericstandalone_i2c_status1 = builder_xilinxmultiregimpl191;
assign main_genericstandalone_i2c_status2 = builder_xilinxmultiregimpl201;
assign main_genericstandalone_rtio_core_sed_lane_dist_enable_spread = builder_xilinxmultiregimpl211;
assign main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_o = builder_xilinxmultiregimpl221;
assign main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_o = builder_xilinxmultiregimpl231;
assign main_genericstandalone_rtio_core_o_collision_sync_data_o = builder_xilinxmultiregimpl241;
assign main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_o = builder_xilinxmultiregimpl251;
assign main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_o = builder_xilinxmultiregimpl261;
assign main_genericstandalone_rtio_core_o_busy_sync_data_o = builder_xilinxmultiregimpl271;
assign main_genericstandalone_mon_bussynchronizer0_o = builder_xilinxmultiregimpl281;
assign main_genericstandalone_mon_bussynchronizer1_o = builder_xilinxmultiregimpl291;
assign main_genericstandalone_mon_bussynchronizer2_o = builder_xilinxmultiregimpl301;
assign main_genericstandalone_mon_bussynchronizer3_o = builder_xilinxmultiregimpl311;
assign main_genericstandalone_mon_bussynchronizer4_o = builder_xilinxmultiregimpl321;
assign main_genericstandalone_mon_bussynchronizer5_o = builder_xilinxmultiregimpl331;
assign main_genericstandalone_mon_bussynchronizer6_o = builder_xilinxmultiregimpl341;
assign main_genericstandalone_mon_bussynchronizer7_o = builder_xilinxmultiregimpl351;
assign main_genericstandalone_mon_bussynchronizer8_o = builder_xilinxmultiregimpl361;
assign main_genericstandalone_mon_bussynchronizer9_o = builder_xilinxmultiregimpl371;
assign main_genericstandalone_mon_bussynchronizer10_o = builder_xilinxmultiregimpl381;
assign main_genericstandalone_mon_bussynchronizer11_o = builder_xilinxmultiregimpl391;
assign main_genericstandalone_mon_bussynchronizer12_o = builder_xilinxmultiregimpl401;
assign main_genericstandalone_mon_bussynchronizer13_o = builder_xilinxmultiregimpl411;
assign main_genericstandalone_mon_bussynchronizer14_o = builder_xilinxmultiregimpl421;
assign main_genericstandalone_mon_bussynchronizer15_o = builder_xilinxmultiregimpl431;
assign main_genericstandalone_mon_bussynchronizer16_o = builder_xilinxmultiregimpl441;
assign main_genericstandalone_mon_bussynchronizer17_o = builder_xilinxmultiregimpl451;
assign main_genericstandalone_mon_bussynchronizer18_o = builder_xilinxmultiregimpl461;
assign main_genericstandalone_mon_bussynchronizer19_o = builder_xilinxmultiregimpl471;
assign main_genericstandalone_mon_bussynchronizer20_ping_toggle_o = builder_xilinxmultiregimpl481;
assign main_genericstandalone_mon_bussynchronizer20_pong_toggle_o = builder_xilinxmultiregimpl491;
assign main_genericstandalone_mon_bussynchronizer20_obuffer = builder_xilinxmultiregimpl501;
assign main_genericstandalone_mon_bussynchronizer21_ping_toggle_o = builder_xilinxmultiregimpl511;
assign main_genericstandalone_mon_bussynchronizer21_pong_toggle_o = builder_xilinxmultiregimpl521;
assign main_genericstandalone_mon_bussynchronizer21_obuffer = builder_xilinxmultiregimpl531;
assign main_genericstandalone_mon_bussynchronizer22_ping_toggle_o = builder_xilinxmultiregimpl541;
assign main_genericstandalone_mon_bussynchronizer22_pong_toggle_o = builder_xilinxmultiregimpl551;
assign main_genericstandalone_mon_bussynchronizer22_obuffer = builder_xilinxmultiregimpl561;
assign main_genericstandalone_mon_bussynchronizer23_ping_toggle_o = builder_xilinxmultiregimpl571;
assign main_genericstandalone_mon_bussynchronizer23_pong_toggle_o = builder_xilinxmultiregimpl581;
assign main_genericstandalone_mon_bussynchronizer23_obuffer = builder_xilinxmultiregimpl591;
assign main_genericstandalone_mon_bussynchronizer24_o = builder_xilinxmultiregimpl601;
assign main_genericstandalone_mon_bussynchronizer25_o = builder_xilinxmultiregimpl611;
assign main_genericstandalone_mon_bussynchronizer26_o = builder_xilinxmultiregimpl621;
assign main_genericstandalone_mon_bussynchronizer27_o = builder_xilinxmultiregimpl631;
assign main_genericstandalone_mon_bussynchronizer28_o = builder_xilinxmultiregimpl641;
assign main_genericstandalone_mon_bussynchronizer29_ping_toggle_o = builder_xilinxmultiregimpl651;
assign main_genericstandalone_mon_bussynchronizer29_pong_toggle_o = builder_xilinxmultiregimpl661;
assign main_genericstandalone_mon_bussynchronizer29_obuffer = builder_xilinxmultiregimpl671;
assign main_genericstandalone_mon_bussynchronizer30_ping_toggle_o = builder_xilinxmultiregimpl681;
assign main_genericstandalone_mon_bussynchronizer30_pong_toggle_o = builder_xilinxmultiregimpl691;
assign main_genericstandalone_mon_bussynchronizer30_obuffer = builder_xilinxmultiregimpl701;
assign main_genericstandalone_mon_bussynchronizer31_ping_toggle_o = builder_xilinxmultiregimpl711;
assign main_genericstandalone_mon_bussynchronizer31_pong_toggle_o = builder_xilinxmultiregimpl721;
assign main_genericstandalone_mon_bussynchronizer31_obuffer = builder_xilinxmultiregimpl731;
assign main_genericstandalone_mon_bussynchronizer32_ping_toggle_o = builder_xilinxmultiregimpl741;
assign main_genericstandalone_mon_bussynchronizer32_pong_toggle_o = builder_xilinxmultiregimpl751;
assign main_genericstandalone_mon_bussynchronizer32_obuffer = builder_xilinxmultiregimpl761;
assign main_genericstandalone_mon_bussynchronizer33_o = builder_xilinxmultiregimpl771;
assign main_genericstandalone_mon_bussynchronizer34_o = builder_xilinxmultiregimpl781;
assign main_genericstandalone_mon_bussynchronizer35_o = builder_xilinxmultiregimpl791;
assign main_genericstandalone_mon_bussynchronizer36_o = builder_xilinxmultiregimpl801;
assign main_genericstandalone_mon_bussynchronizer37_o = builder_xilinxmultiregimpl811;
assign main_genericstandalone_mon_bussynchronizer38_o = builder_xilinxmultiregimpl821;
assign main_genericstandalone_mon_bussynchronizer39_ping_toggle_o = builder_xilinxmultiregimpl831;
assign main_genericstandalone_mon_bussynchronizer39_pong_toggle_o = builder_xilinxmultiregimpl841;
assign main_genericstandalone_mon_bussynchronizer39_obuffer = builder_xilinxmultiregimpl851;
assign main_genericstandalone_mon_bussynchronizer40_ping_toggle_o = builder_xilinxmultiregimpl861;
assign main_genericstandalone_mon_bussynchronizer40_pong_toggle_o = builder_xilinxmultiregimpl871;
assign main_genericstandalone_mon_bussynchronizer40_obuffer = builder_xilinxmultiregimpl881;
assign main_genericstandalone_mon_bussynchronizer41_ping_toggle_o = builder_xilinxmultiregimpl891;
assign main_genericstandalone_mon_bussynchronizer41_pong_toggle_o = builder_xilinxmultiregimpl901;
assign main_genericstandalone_mon_bussynchronizer41_obuffer = builder_xilinxmultiregimpl911;
assign main_genericstandalone_mon_bussynchronizer42_ping_toggle_o = builder_xilinxmultiregimpl921;
assign main_genericstandalone_mon_bussynchronizer42_pong_toggle_o = builder_xilinxmultiregimpl931;
assign main_genericstandalone_mon_bussynchronizer42_obuffer = builder_xilinxmultiregimpl941;
assign main_genericstandalone_mon_bussynchronizer43_ping_toggle_o = builder_xilinxmultiregimpl951;
assign main_genericstandalone_mon_bussynchronizer43_pong_toggle_o = builder_xilinxmultiregimpl961;
assign main_genericstandalone_mon_bussynchronizer43_obuffer = builder_xilinxmultiregimpl971;
assign main_genericstandalone_mon_bussynchronizer44_ping_toggle_o = builder_xilinxmultiregimpl981;
assign main_genericstandalone_mon_bussynchronizer44_pong_toggle_o = builder_xilinxmultiregimpl991;
assign main_genericstandalone_mon_bussynchronizer44_obuffer = builder_xilinxmultiregimpl1001;
assign main_genericstandalone_mon_bussynchronizer45_ping_toggle_o = builder_xilinxmultiregimpl1011;
assign main_genericstandalone_mon_bussynchronizer45_pong_toggle_o = builder_xilinxmultiregimpl1021;
assign main_genericstandalone_mon_bussynchronizer45_obuffer = builder_xilinxmultiregimpl1031;
assign main_genericstandalone_mon_bussynchronizer46_ping_toggle_o = builder_xilinxmultiregimpl1041;
assign main_genericstandalone_mon_bussynchronizer46_pong_toggle_o = builder_xilinxmultiregimpl1051;
assign main_genericstandalone_mon_bussynchronizer46_obuffer = builder_xilinxmultiregimpl1061;
assign main_genericstandalone_mon_bussynchronizer47_ping_toggle_o = builder_xilinxmultiregimpl1071;
assign main_genericstandalone_mon_bussynchronizer47_pong_toggle_o = builder_xilinxmultiregimpl1081;
assign main_genericstandalone_mon_bussynchronizer47_obuffer = builder_xilinxmultiregimpl1091;
assign main_genericstandalone_mon_bussynchronizer48_ping_toggle_o = builder_xilinxmultiregimpl1101;
assign main_genericstandalone_mon_bussynchronizer48_pong_toggle_o = builder_xilinxmultiregimpl1111;
assign main_genericstandalone_mon_bussynchronizer48_obuffer = builder_xilinxmultiregimpl1121;
assign main_genericstandalone_mon_bussynchronizer49_ping_toggle_o = builder_xilinxmultiregimpl1131;
assign main_genericstandalone_mon_bussynchronizer49_pong_toggle_o = builder_xilinxmultiregimpl1141;
assign main_genericstandalone_mon_bussynchronizer49_obuffer = builder_xilinxmultiregimpl1151;
assign main_genericstandalone_mon_bussynchronizer50_ping_toggle_o = builder_xilinxmultiregimpl1161;
assign main_genericstandalone_mon_bussynchronizer50_pong_toggle_o = builder_xilinxmultiregimpl1171;
assign main_genericstandalone_mon_bussynchronizer50_obuffer = builder_xilinxmultiregimpl1181;
assign main_genericstandalone_mon_bussynchronizer51_ping_toggle_o = builder_xilinxmultiregimpl1191;
assign main_genericstandalone_mon_bussynchronizer51_pong_toggle_o = builder_xilinxmultiregimpl1201;
assign main_genericstandalone_mon_bussynchronizer51_obuffer = builder_xilinxmultiregimpl1211;
assign main_genericstandalone_mon_bussynchronizer52_ping_toggle_o = builder_xilinxmultiregimpl1221;
assign main_genericstandalone_mon_bussynchronizer52_pong_toggle_o = builder_xilinxmultiregimpl1231;
assign main_genericstandalone_mon_bussynchronizer52_obuffer = builder_xilinxmultiregimpl1241;
assign main_genericstandalone_mon_bussynchronizer53_ping_toggle_o = builder_xilinxmultiregimpl1251;
assign main_genericstandalone_mon_bussynchronizer53_pong_toggle_o = builder_xilinxmultiregimpl1261;
assign main_genericstandalone_mon_bussynchronizer53_obuffer = builder_xilinxmultiregimpl1271;
assign main_genericstandalone_mon_bussynchronizer54_ping_toggle_o = builder_xilinxmultiregimpl1281;
assign main_genericstandalone_mon_bussynchronizer54_pong_toggle_o = builder_xilinxmultiregimpl1291;
assign main_genericstandalone_mon_bussynchronizer54_obuffer = builder_xilinxmultiregimpl1301;
assign main_genericstandalone_mon_bussynchronizer55_ping_toggle_o = builder_xilinxmultiregimpl1311;
assign main_genericstandalone_mon_bussynchronizer55_pong_toggle_o = builder_xilinxmultiregimpl1321;
assign main_genericstandalone_mon_bussynchronizer55_obuffer = builder_xilinxmultiregimpl1331;
assign main_genericstandalone_mon_bussynchronizer56_ping_toggle_o = builder_xilinxmultiregimpl1341;
assign main_genericstandalone_mon_bussynchronizer56_pong_toggle_o = builder_xilinxmultiregimpl1351;
assign main_genericstandalone_mon_bussynchronizer56_obuffer = builder_xilinxmultiregimpl1361;
assign main_genericstandalone_mon_bussynchronizer57_ping_toggle_o = builder_xilinxmultiregimpl1371;
assign main_genericstandalone_mon_bussynchronizer57_pong_toggle_o = builder_xilinxmultiregimpl1381;
assign main_genericstandalone_mon_bussynchronizer57_obuffer = builder_xilinxmultiregimpl1391;
assign main_genericstandalone_mon_bussynchronizer58_ping_toggle_o = builder_xilinxmultiregimpl1401;
assign main_genericstandalone_mon_bussynchronizer58_pong_toggle_o = builder_xilinxmultiregimpl1411;
assign main_genericstandalone_mon_bussynchronizer58_obuffer = builder_xilinxmultiregimpl1421;
assign main_genericstandalone_mon_bussynchronizer59_ping_toggle_o = builder_xilinxmultiregimpl1431;
assign main_genericstandalone_mon_bussynchronizer59_pong_toggle_o = builder_xilinxmultiregimpl1441;
assign main_genericstandalone_mon_bussynchronizer59_obuffer = builder_xilinxmultiregimpl1451;
assign main_genericstandalone_mon_bussynchronizer60_ping_toggle_o = builder_xilinxmultiregimpl1461;
assign main_genericstandalone_mon_bussynchronizer60_pong_toggle_o = builder_xilinxmultiregimpl1471;
assign main_genericstandalone_mon_bussynchronizer60_obuffer = builder_xilinxmultiregimpl1481;
assign main_genericstandalone_mon_bussynchronizer61_ping_toggle_o = builder_xilinxmultiregimpl1491;
assign main_genericstandalone_mon_bussynchronizer61_pong_toggle_o = builder_xilinxmultiregimpl1501;
assign main_genericstandalone_mon_bussynchronizer61_obuffer = builder_xilinxmultiregimpl1511;
assign main_genericstandalone_mon_bussynchronizer62_ping_toggle_o = builder_xilinxmultiregimpl1521;
assign main_genericstandalone_mon_bussynchronizer62_pong_toggle_o = builder_xilinxmultiregimpl1531;
assign main_genericstandalone_mon_bussynchronizer62_obuffer = builder_xilinxmultiregimpl1541;
assign main_genericstandalone_mon_bussynchronizer63_ping_toggle_o = builder_xilinxmultiregimpl1551;
assign main_genericstandalone_mon_bussynchronizer63_pong_toggle_o = builder_xilinxmultiregimpl1561;
assign main_genericstandalone_mon_bussynchronizer63_obuffer = builder_xilinxmultiregimpl1571;
assign main_genericstandalone_mon_bussynchronizer64_ping_toggle_o = builder_xilinxmultiregimpl1581;
assign main_genericstandalone_mon_bussynchronizer64_pong_toggle_o = builder_xilinxmultiregimpl1591;
assign main_genericstandalone_mon_bussynchronizer64_obuffer = builder_xilinxmultiregimpl1601;
assign main_genericstandalone_mon_bussynchronizer65_ping_toggle_o = builder_xilinxmultiregimpl1611;
assign main_genericstandalone_mon_bussynchronizer65_pong_toggle_o = builder_xilinxmultiregimpl1621;
assign main_genericstandalone_mon_bussynchronizer65_obuffer = builder_xilinxmultiregimpl1631;
assign main_genericstandalone_mon_bussynchronizer66_ping_toggle_o = builder_xilinxmultiregimpl1641;
assign main_genericstandalone_mon_bussynchronizer66_pong_toggle_o = builder_xilinxmultiregimpl1651;
assign main_genericstandalone_mon_bussynchronizer66_obuffer = builder_xilinxmultiregimpl1661;
assign main_genericstandalone_mon_bussynchronizer67_ping_toggle_o = builder_xilinxmultiregimpl1671;
assign main_genericstandalone_mon_bussynchronizer67_pong_toggle_o = builder_xilinxmultiregimpl1681;
assign main_genericstandalone_mon_bussynchronizer67_obuffer = builder_xilinxmultiregimpl1691;
assign main_genericstandalone_mon_bussynchronizer68_ping_toggle_o = builder_xilinxmultiregimpl1701;
assign main_genericstandalone_mon_bussynchronizer68_pong_toggle_o = builder_xilinxmultiregimpl1711;
assign main_genericstandalone_mon_bussynchronizer68_obuffer = builder_xilinxmultiregimpl1721;
assign main_genericstandalone_mon_bussynchronizer69_ping_toggle_o = builder_xilinxmultiregimpl1731;
assign main_genericstandalone_mon_bussynchronizer69_pong_toggle_o = builder_xilinxmultiregimpl1741;
assign main_genericstandalone_mon_bussynchronizer69_obuffer = builder_xilinxmultiregimpl1751;
assign main_genericstandalone_mon_bussynchronizer70_ping_toggle_o = builder_xilinxmultiregimpl1761;
assign main_genericstandalone_mon_bussynchronizer70_pong_toggle_o = builder_xilinxmultiregimpl1771;
assign main_genericstandalone_mon_bussynchronizer70_obuffer = builder_xilinxmultiregimpl1781;
assign main_genericstandalone_mon_bussynchronizer71_o = builder_xilinxmultiregimpl1791;
assign main_genericstandalone_mon_bussynchronizer72_o = builder_xilinxmultiregimpl1801;
assign main_genericstandalone_mon_bussynchronizer73_o = builder_xilinxmultiregimpl1811;
assign main_genericstandalone_mon_bussynchronizer74_o = builder_xilinxmultiregimpl1821;
assign main_genericstandalone_mon_bussynchronizer75_o = builder_xilinxmultiregimpl1831;
assign main_inout_8x0_inout_8x0_override_en = builder_xilinxmultiregimpl1841;
assign main_inout_8x0_inout_8x0_override_o = builder_xilinxmultiregimpl1851;
assign main_inout_8x0_inout_8x0_override_oe = builder_xilinxmultiregimpl1861;
assign main_inout_8x1_inout_8x1_override_en = builder_xilinxmultiregimpl1871;
assign main_inout_8x1_inout_8x1_override_o = builder_xilinxmultiregimpl1881;
assign main_inout_8x1_inout_8x1_override_oe = builder_xilinxmultiregimpl1891;
assign main_inout_8x2_inout_8x2_override_en = builder_xilinxmultiregimpl1901;
assign main_inout_8x2_inout_8x2_override_o = builder_xilinxmultiregimpl1911;
assign main_inout_8x2_inout_8x2_override_oe = builder_xilinxmultiregimpl1921;
assign main_inout_8x3_inout_8x3_override_en = builder_xilinxmultiregimpl1931;
assign main_inout_8x3_inout_8x3_override_o = builder_xilinxmultiregimpl1941;
assign main_inout_8x3_inout_8x3_override_oe = builder_xilinxmultiregimpl1951;
assign main_output_8x0_override_en0 = builder_xilinxmultiregimpl1961;
assign main_output_8x0_override_o0 = builder_xilinxmultiregimpl1971;
assign main_output_8x1_override_en0 = builder_xilinxmultiregimpl1981;
assign main_output_8x1_override_o0 = builder_xilinxmultiregimpl1991;
assign main_output_8x2_override_en = builder_xilinxmultiregimpl2001;
assign main_output_8x2_override_o = builder_xilinxmultiregimpl2011;
assign main_output_8x3_override_en = builder_xilinxmultiregimpl2021;
assign main_output_8x3_override_o = builder_xilinxmultiregimpl2031;
assign main_output_8x4_override_en = builder_xilinxmultiregimpl2041;
assign main_output_8x4_override_o = builder_xilinxmultiregimpl2051;
assign main_output_8x5_override_en = builder_xilinxmultiregimpl2061;
assign main_output_8x5_override_o = builder_xilinxmultiregimpl2071;
assign main_output_8x6_override_en = builder_xilinxmultiregimpl2081;
assign main_output_8x6_override_o = builder_xilinxmultiregimpl2091;
assign main_output_8x7_override_en = builder_xilinxmultiregimpl2101;
assign main_output_8x7_override_o = builder_xilinxmultiregimpl2111;
assign main_output_8x8_override_en = builder_xilinxmultiregimpl2121;
assign main_output_8x8_override_o = builder_xilinxmultiregimpl2131;
assign main_output_8x9_override_en = builder_xilinxmultiregimpl2141;
assign main_output_8x9_override_o = builder_xilinxmultiregimpl2151;
assign main_output_8x10_override_en = builder_xilinxmultiregimpl2161;
assign main_output_8x10_override_o = builder_xilinxmultiregimpl2171;
assign main_output_8x11_override_en = builder_xilinxmultiregimpl2181;
assign main_output_8x11_override_o = builder_xilinxmultiregimpl2191;
assign main_output_8x0_override_en1 = builder_xilinxmultiregimpl2201;
assign main_output_8x0_override_o1 = builder_xilinxmultiregimpl2211;
assign main_output_8x12_override_en = builder_xilinxmultiregimpl2221;
assign main_output_8x12_override_o = builder_xilinxmultiregimpl2231;
assign main_output_8x13_override_en = builder_xilinxmultiregimpl2241;
assign main_output_8x13_override_o = builder_xilinxmultiregimpl2251;
assign main_output_8x14_override_en = builder_xilinxmultiregimpl2261;
assign main_output_8x14_override_o = builder_xilinxmultiregimpl2271;
assign main_output_8x15_override_en = builder_xilinxmultiregimpl2281;
assign main_output_8x15_override_o = builder_xilinxmultiregimpl2291;
assign main_output_8x1_override_en1 = builder_xilinxmultiregimpl2301;
assign main_output_8x1_override_o1 = builder_xilinxmultiregimpl2311;
assign main_output_8x16_override_en = builder_xilinxmultiregimpl2321;
assign main_output_8x16_override_o = builder_xilinxmultiregimpl2331;
assign main_output_8x17_override_en = builder_xilinxmultiregimpl2341;
assign main_output_8x17_override_o = builder_xilinxmultiregimpl2351;
assign main_output_8x18_override_en = builder_xilinxmultiregimpl2361;
assign main_output_8x18_override_o = builder_xilinxmultiregimpl2371;
assign main_output_8x19_override_en = builder_xilinxmultiregimpl2381;
assign main_output_8x19_override_o = builder_xilinxmultiregimpl2391;
assign main_output_8x20_override_en = builder_xilinxmultiregimpl2401;
assign main_output_8x20_override_o = builder_xilinxmultiregimpl2411;
assign main_ldac_phy_override_en = builder_xilinxmultiregimpl2421;
assign main_ldac_phy_override_o = builder_xilinxmultiregimpl2431;
assign main_clr_phy_override_en = builder_xilinxmultiregimpl2441;
assign main_clr_phy_override_o = builder_xilinxmultiregimpl2451;
assign main_output0_override_en = builder_xilinxmultiregimpl2461;
assign main_output0_override_o = builder_xilinxmultiregimpl2471;
assign main_output1_override_en = builder_xilinxmultiregimpl2481;
assign main_output1_override_o = builder_xilinxmultiregimpl2491;
assign main_output2_override_en = builder_xilinxmultiregimpl2501;
assign main_output2_override_o = builder_xilinxmultiregimpl2511;

always @(posedge bootstrap_clk) begin
	main_genericstandalone_genericstandalone_crg_o_clk_sw <= main_genericstandalone_genericstandalone_crg_o_switch;
	main_genericstandalone_genericstandalone_crg_o_reset <= main_genericstandalone_genericstandalone_crg_reset;
	builder_rtiosyscrg_state <= builder_rtiosyscrg_next_state;
	if (main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value_ce0) begin
		main_genericstandalone_genericstandalone_crg_delay_counter <= main_genericstandalone_genericstandalone_crg_delay_counter_rtiosyscrg_next_value0;
	end
	if (main_genericstandalone_genericstandalone_crg_o_switch_rtiosyscrg_next_value_ce1) begin
		main_genericstandalone_genericstandalone_crg_o_switch <= main_genericstandalone_genericstandalone_crg_o_switch_rtiosyscrg_next_value1;
	end
	builder_xilinxmultiregimpl10 <= main_genericstandalone_genericstandalone_crg_i_clk_sw;
	builder_xilinxmultiregimpl11 <= builder_xilinxmultiregimpl10;
end

always @(posedge clk200_clk) begin
	if ((main_genericstandalone_genericstandalone_crg_reset_counter != 1'd0)) begin
		main_genericstandalone_genericstandalone_crg_reset_counter <= (main_genericstandalone_genericstandalone_crg_reset_counter - 1'd1);
	end else begin
		main_genericstandalone_genericstandalone_crg_ic_reset <= 1'd0;
	end
	if (clk200_rst) begin
		main_genericstandalone_genericstandalone_crg_reset_counter <= 4'd15;
		main_genericstandalone_genericstandalone_crg_ic_reset <= 1'd1;
	end
end

always @(posedge eth_rx_clk) begin
	main_genericstandalone_pcs_rx_en_d <= main_genericstandalone_pcs_receivepath_rx_en;
	main_genericstandalone_pcs_source_stb <= main_genericstandalone_pcs_receivepath_sample_en;
	main_genericstandalone_pcs_source_payload_data <= main_genericstandalone_pcs_receivepath_rx_data;
	if (main_genericstandalone_pcs_receivepath_seen_config_reg) begin
		main_genericstandalone_pcs_c_counter <= 3'd4;
	end else begin
		if ((main_genericstandalone_pcs_c_counter != 1'd0)) begin
			main_genericstandalone_pcs_c_counter <= (main_genericstandalone_pcs_c_counter - 1'd1);
		end
	end
	main_genericstandalone_pcs_rx_config_reg_abi_i <= 1'd0;
	main_genericstandalone_pcs_rx_config_reg_ack_i <= 1'd0;
	if (main_genericstandalone_pcs_receivepath_seen_config_reg) begin
		main_genericstandalone_pcs_prev_config_reg <= main_genericstandalone_pcs_receivepath_config_reg;
		if (((main_genericstandalone_pcs_c_counter == 1'd1) & ((main_genericstandalone_pcs_prev_config_reg & 16'd49151) == (main_genericstandalone_pcs_receivepath_config_reg & 16'd49151)))) begin
			if ((main_genericstandalone_pcs_prev_config_reg[14] & main_genericstandalone_pcs_receivepath_config_reg[14])) begin
				main_genericstandalone_pcs_rx_config_reg_ack_i <= 1'd1;
			end else begin
				main_genericstandalone_pcs_rx_config_reg_abi_i <= 1'd1;
			end
		end
		main_genericstandalone_pcs_lp_abi_i <= main_genericstandalone_pcs_receivepath_config_reg;
	end
	main_genericstandalone_pcs_receivepath_seen_config_reg <= 1'd0;
	if (main_genericstandalone_pcs_receivepath_load_config_reg_lsb) begin
		main_genericstandalone_pcs_receivepath_config_reg_lsb <= main_genericstandalone_pcs_receivepath_d;
	end
	if (main_genericstandalone_pcs_receivepath_load_config_reg_msb) begin
		main_genericstandalone_pcs_receivepath_config_reg <= {main_genericstandalone_pcs_receivepath_d, main_genericstandalone_pcs_receivepath_config_reg_lsb};
		main_genericstandalone_pcs_receivepath_seen_config_reg <= 1'd1;
	end
	if (((~main_genericstandalone_pcs_receivepath_timer_en) | (main_genericstandalone_pcs_receivepath_timer == 1'd0))) begin
		if ((main_genericstandalone_pcs_receivepath_sgmii_speed == 1'd0)) begin
			main_genericstandalone_pcs_receivepath_timer <= 7'd99;
		end else begin
			if ((main_genericstandalone_pcs_receivepath_sgmii_speed == 1'd1)) begin
				main_genericstandalone_pcs_receivepath_timer <= 4'd9;
			end else begin
				if ((main_genericstandalone_pcs_receivepath_sgmii_speed == 2'd2)) begin
					main_genericstandalone_pcs_receivepath_timer <= 1'd0;
				end
			end
		end
	end else begin
		if (main_genericstandalone_pcs_receivepath_timer_en) begin
			main_genericstandalone_pcs_receivepath_timer <= (main_genericstandalone_pcs_receivepath_timer - 1'd1);
		end
	end
	main_genericstandalone_pcs_receivepath_k <= 1'd0;
	if ((main_genericstandalone_pcs_receivepath_input_msb_first[9:4] == 4'd15)) begin
		main_genericstandalone_pcs_receivepath_k <= 1'd1;
		main_genericstandalone_pcs_receivepath_code3b <= builder_sync_t_rhs_self0;
	end else begin
		if ((main_genericstandalone_pcs_receivepath_input_msb_first[9:4] == 6'd48)) begin
			main_genericstandalone_pcs_receivepath_k <= 1'd1;
			main_genericstandalone_pcs_receivepath_code3b <= builder_sync_f_t_self0;
		end else begin
			if (((main_genericstandalone_pcs_receivepath_input_msb_first[3:0] == 3'd7) | (main_genericstandalone_pcs_receivepath_input_msb_first[3:0] == 4'd8))) begin
				if (((((((main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 6'd35) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 5'd19)) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 4'd11)) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 6'd52)) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 6'd44)) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 5'd28))) begin
					main_genericstandalone_pcs_receivepath_k <= 1'd1;
				end
			end
			main_genericstandalone_pcs_receivepath_code3b <= builder_sync_f_rhs_self0;
		end
	end
	main_genericstandalone_pcs_receivepath_code5b <= builder_sync_rhs_self0;
	builder_a7_1000basex_receivepath_state <= builder_a7_1000basex_receivepath_next_state;
	main_genericstandalone_pcs_lp_abi_starter <= 1'd0;
	if (main_genericstandalone_pcs_lp_abi_pong_o) begin
		main_genericstandalone_pcs_lp_abi_ibuffer <= main_genericstandalone_pcs_lp_abi_i;
	end
	if (main_genericstandalone_pcs_lp_abi_ping_i) begin
		main_genericstandalone_pcs_lp_abi_ping_toggle_i <= (~main_genericstandalone_pcs_lp_abi_ping_toggle_i);
	end
	main_genericstandalone_pcs_lp_abi_pong_toggle_o_r <= main_genericstandalone_pcs_lp_abi_pong_toggle_o;
	if (main_genericstandalone_pcs_lp_abi_wait) begin
		if ((~main_genericstandalone_pcs_lp_abi_done)) begin
			main_genericstandalone_pcs_lp_abi_count <= (main_genericstandalone_pcs_lp_abi_count - 1'd1);
		end
	end else begin
		main_genericstandalone_pcs_lp_abi_count <= 8'd128;
	end
	if (main_genericstandalone_pcs_seen_valid_ci_i) begin
		main_genericstandalone_pcs_seen_valid_ci_toggle_i <= (~main_genericstandalone_pcs_seen_valid_ci_toggle_i);
	end
	if (main_genericstandalone_pcs_rx_config_reg_abi_i) begin
		main_genericstandalone_pcs_rx_config_reg_abi_toggle_i <= (~main_genericstandalone_pcs_rx_config_reg_abi_toggle_i);
	end
	if (main_genericstandalone_pcs_rx_config_reg_ack_i) begin
		main_genericstandalone_pcs_rx_config_reg_ack_toggle_i <= (~main_genericstandalone_pcs_rx_config_reg_ack_toggle_i);
	end
	if ((main_genericstandalone_phase_half == main_genericstandalone_phase_half_rereg)) begin
		main_genericstandalone_rx_data1 <= main_genericstandalone_rx_data_half[19:10];
	end else begin
		main_genericstandalone_rx_data1 <= main_genericstandalone_rx_data_half[9:0];
	end
	main_genericstandalone_phase_half <= (~main_genericstandalone_phase_half);
	builder_liteethmacpreamblechecker_state <= builder_liteethmacpreamblechecker_next_state;
	if (main_genericstandalone_crc32_checker_crc_ce) begin
		main_genericstandalone_crc32_checker_crc_reg <= main_genericstandalone_crc32_checker_crc_next;
	end
	if (main_genericstandalone_crc32_checker_crc_reset) begin
		main_genericstandalone_crc32_checker_crc_reg <= 32'd4294967295;
	end
	if (((main_genericstandalone_crc32_checker_syncfifo_syncfifo_we & main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable) & (~main_genericstandalone_crc32_checker_syncfifo_replace))) begin
		if ((main_genericstandalone_crc32_checker_syncfifo_produce == 3'd4)) begin
			main_genericstandalone_crc32_checker_syncfifo_produce <= 1'd0;
		end else begin
			main_genericstandalone_crc32_checker_syncfifo_produce <= (main_genericstandalone_crc32_checker_syncfifo_produce + 1'd1);
		end
	end
	if (main_genericstandalone_crc32_checker_syncfifo_do_read) begin
		if ((main_genericstandalone_crc32_checker_syncfifo_consume == 3'd4)) begin
			main_genericstandalone_crc32_checker_syncfifo_consume <= 1'd0;
		end else begin
			main_genericstandalone_crc32_checker_syncfifo_consume <= (main_genericstandalone_crc32_checker_syncfifo_consume + 1'd1);
		end
	end
	if (((main_genericstandalone_crc32_checker_syncfifo_syncfifo_we & main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable) & (~main_genericstandalone_crc32_checker_syncfifo_replace))) begin
		if ((~main_genericstandalone_crc32_checker_syncfifo_do_read)) begin
			main_genericstandalone_crc32_checker_syncfifo_level <= (main_genericstandalone_crc32_checker_syncfifo_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_crc32_checker_syncfifo_do_read) begin
			main_genericstandalone_crc32_checker_syncfifo_level <= (main_genericstandalone_crc32_checker_syncfifo_level - 1'd1);
		end
	end
	if (main_genericstandalone_crc32_checker_fifo_reset) begin
		main_genericstandalone_crc32_checker_syncfifo_level <= 3'd0;
		main_genericstandalone_crc32_checker_syncfifo_produce <= 3'd0;
		main_genericstandalone_crc32_checker_syncfifo_consume <= 3'd0;
	end
	builder_liteethmaccrc32checker_state <= builder_liteethmaccrc32checker_next_state;
	if (main_genericstandalone_ps_preamble_error_i) begin
		main_genericstandalone_ps_preamble_error_toggle_i <= (~main_genericstandalone_ps_preamble_error_toggle_i);
	end
	if (main_genericstandalone_ps_crc_error_i) begin
		main_genericstandalone_ps_crc_error_toggle_i <= (~main_genericstandalone_ps_crc_error_toggle_i);
	end
	if (main_genericstandalone_rx_converter_converter_source_ack) begin
		main_genericstandalone_rx_converter_converter_strobe_all <= 1'd0;
	end
	if (main_genericstandalone_rx_converter_converter_load_part) begin
		if (((main_genericstandalone_rx_converter_converter_demux == 3'd7) | main_genericstandalone_rx_converter_converter_sink_eop)) begin
			main_genericstandalone_rx_converter_converter_demux <= 1'd0;
			main_genericstandalone_rx_converter_converter_strobe_all <= 1'd1;
		end else begin
			main_genericstandalone_rx_converter_converter_demux <= (main_genericstandalone_rx_converter_converter_demux + 1'd1);
		end
	end
	if ((main_genericstandalone_rx_converter_converter_source_stb & main_genericstandalone_rx_converter_converter_source_ack)) begin
		main_genericstandalone_rx_converter_converter_source_eop <= main_genericstandalone_rx_converter_converter_sink_eop;
	end else begin
		if ((main_genericstandalone_rx_converter_converter_sink_stb & main_genericstandalone_rx_converter_converter_sink_ack)) begin
			main_genericstandalone_rx_converter_converter_source_eop <= (main_genericstandalone_rx_converter_converter_sink_eop | main_genericstandalone_rx_converter_converter_source_eop);
		end
	end
	if (main_genericstandalone_rx_converter_converter_load_part) begin
		case (main_genericstandalone_rx_converter_converter_demux)
			1'd0: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[9:0] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			1'd1: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[19:10] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			2'd2: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[29:20] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			2'd3: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[39:30] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			3'd4: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[49:40] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			3'd5: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[59:50] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			3'd6: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[69:60] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			3'd7: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[79:70] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
		endcase
	end
	main_genericstandalone_rx_cdc_graycounter0_q_binary <= main_genericstandalone_rx_cdc_graycounter0_q_next_binary;
	main_genericstandalone_rx_cdc_graycounter0_q <= main_genericstandalone_rx_cdc_graycounter0_q_next;
	if (eth_rx_rst) begin
		main_genericstandalone_pcs_receivepath_seen_config_reg <= 1'd0;
		main_genericstandalone_pcs_receivepath_config_reg <= 16'd0;
		main_genericstandalone_pcs_receivepath_k <= 1'd0;
		main_genericstandalone_pcs_receivepath_code5b <= 5'd0;
		main_genericstandalone_pcs_receivepath_code3b <= 3'd0;
		main_genericstandalone_pcs_receivepath_config_reg_lsb <= 8'd0;
		main_genericstandalone_pcs_receivepath_timer <= 10'd0;
		main_genericstandalone_pcs_source_stb <= 1'd0;
		main_genericstandalone_pcs_source_payload_data <= 8'd0;
		main_genericstandalone_pcs_lp_abi_i <= 16'd0;
		main_genericstandalone_pcs_lp_abi_starter <= 1'd1;
		main_genericstandalone_pcs_lp_abi_count <= 8'd128;
		main_genericstandalone_pcs_rx_en_d <= 1'd0;
		main_genericstandalone_pcs_rx_config_reg_abi_i <= 1'd0;
		main_genericstandalone_pcs_rx_config_reg_ack_i <= 1'd0;
		main_genericstandalone_pcs_c_counter <= 3'd0;
		main_genericstandalone_pcs_prev_config_reg <= 16'd0;
		main_genericstandalone_rx_data1 <= 10'd0;
		main_genericstandalone_phase_half <= 1'd0;
		main_genericstandalone_crc32_checker_crc_reg <= 32'd4294967295;
		main_genericstandalone_crc32_checker_syncfifo_level <= 3'd0;
		main_genericstandalone_crc32_checker_syncfifo_produce <= 3'd0;
		main_genericstandalone_crc32_checker_syncfifo_consume <= 3'd0;
		main_genericstandalone_rx_converter_converter_source_eop <= 1'd0;
		main_genericstandalone_rx_converter_converter_source_payload_data <= 80'd0;
		main_genericstandalone_rx_converter_converter_demux <= 3'd0;
		main_genericstandalone_rx_converter_converter_strobe_all <= 1'd0;
		main_genericstandalone_rx_cdc_graycounter0_q <= 7'd0;
		main_genericstandalone_rx_cdc_graycounter0_q_binary <= 7'd0;
		builder_a7_1000basex_receivepath_state <= 3'd0;
		builder_liteethmacpreamblechecker_state <= 1'd0;
		builder_liteethmaccrc32checker_state <= 2'd0;
	end
	builder_xilinxmultiregimpl50 <= main_genericstandalone_pcs_lp_abi_pong_toggle_i;
	builder_xilinxmultiregimpl51 <= builder_xilinxmultiregimpl50;
	builder_xilinxmultiregimpl180 <= main_genericstandalone_rx_cdc_graycounter1_q;
	builder_xilinxmultiregimpl181 <= builder_xilinxmultiregimpl180;
end

always @(posedge eth_rx_half_clk) begin
	main_genericstandalone_phase_half_rereg <= main_genericstandalone_phase_half;
end

always @(posedge eth_tx_clk) begin
	main_genericstandalone_pcs_checker_tick <= 1'd0;
	if ((main_genericstandalone_pcs_checker_counter == 1'd0)) begin
		main_genericstandalone_pcs_checker_tick <= 1'd1;
		main_genericstandalone_pcs_checker_counter <= 20'd750000;
	end else begin
		main_genericstandalone_pcs_checker_counter <= (main_genericstandalone_pcs_checker_counter - 1'd1);
	end
	if (main_genericstandalone_pcs_seen_valid_ci_o) begin
		main_genericstandalone_pcs_checker_ok <= 1'd1;
	end
	if (main_genericstandalone_pcs_checker_tick) begin
		main_genericstandalone_pcs_checker_ok <= 1'd0;
	end
	main_genericstandalone_pcs_transmitpath_parity <= (~main_genericstandalone_pcs_transmitpath_parity);
	if (main_genericstandalone_pcs_transmitpath_load_config_reg_buffer) begin
		main_genericstandalone_pcs_transmitpath_config_reg_buffer <= main_genericstandalone_pcs_transmitpath_config_reg;
	end
	if (((~main_genericstandalone_pcs_transmitpath_timer_en) | (main_genericstandalone_pcs_transmitpath_timer == 1'd0))) begin
		if ((main_genericstandalone_pcs_transmitpath_sgmii_speed == 1'd0)) begin
			main_genericstandalone_pcs_transmitpath_timer <= 7'd99;
		end else begin
			if ((main_genericstandalone_pcs_transmitpath_sgmii_speed == 1'd1)) begin
				main_genericstandalone_pcs_transmitpath_timer <= 4'd9;
			end else begin
				if ((main_genericstandalone_pcs_transmitpath_sgmii_speed == 2'd2)) begin
					main_genericstandalone_pcs_transmitpath_timer <= 1'd0;
				end
			end
		end
	end else begin
		if (main_genericstandalone_pcs_transmitpath_timer_en) begin
			main_genericstandalone_pcs_transmitpath_timer <= (main_genericstandalone_pcs_transmitpath_timer - 1'd1);
		end
	end
	main_genericstandalone_pcs_transmitpath_encoder_disp_in <= main_genericstandalone_pcs_transmitpath_encoder_disp_out;
	main_genericstandalone_pcs_transmitpath_encoder2 <= main_genericstandalone_pcs_transmitpath_encoder_output;
	main_genericstandalone_pcs_transmitpath_encoder3 <= main_genericstandalone_pcs_transmitpath_encoder_disp_out;
	if ((main_genericstandalone_pcs_transmitpath_encoder_k & (main_genericstandalone_pcs_transmitpath_encoder_d[4:0] == 5'd28))) begin
		main_genericstandalone_pcs_transmitpath_encoder_code6b <= 6'd48;
		main_genericstandalone_pcs_transmitpath_encoder_code6b_unbalanced <= 1'd1;
		main_genericstandalone_pcs_transmitpath_encoder_code6b_flip <= 1'd1;
	end else begin
		main_genericstandalone_pcs_transmitpath_encoder_code6b <= builder_sync_f_rhs_self1;
		main_genericstandalone_pcs_transmitpath_encoder_code6b_unbalanced <= builder_sync_f_rhs_self2;
		main_genericstandalone_pcs_transmitpath_encoder_code6b_flip <= builder_sync_f_rhs_self3;
	end
	main_genericstandalone_pcs_transmitpath_encoder_code4b <= builder_sync_rhs_self1;
	main_genericstandalone_pcs_transmitpath_encoder_code4b_unbalanced <= builder_sync_rhs_self2;
	if (main_genericstandalone_pcs_transmitpath_encoder_k) begin
		main_genericstandalone_pcs_transmitpath_encoder_code4b_flip <= 1'd1;
	end else begin
		main_genericstandalone_pcs_transmitpath_encoder_code4b_flip <= builder_sync_f_rhs_self4;
	end
	main_genericstandalone_pcs_transmitpath_encoder_alt7_rd0 <= 1'd0;
	main_genericstandalone_pcs_transmitpath_encoder_alt7_rd1 <= 1'd0;
	if ((main_genericstandalone_pcs_transmitpath_encoder_d[7:5] == 3'd7)) begin
		if ((((main_genericstandalone_pcs_transmitpath_encoder_d[4:0] == 5'd17) | (main_genericstandalone_pcs_transmitpath_encoder_d[4:0] == 5'd18)) | (main_genericstandalone_pcs_transmitpath_encoder_d[4:0] == 5'd20))) begin
			main_genericstandalone_pcs_transmitpath_encoder_alt7_rd0 <= 1'd1;
		end
		if ((((main_genericstandalone_pcs_transmitpath_encoder_d[4:0] == 4'd11) | (main_genericstandalone_pcs_transmitpath_encoder_d[4:0] == 4'd13)) | (main_genericstandalone_pcs_transmitpath_encoder_d[4:0] == 4'd14))) begin
			main_genericstandalone_pcs_transmitpath_encoder_alt7_rd1 <= 1'd1;
		end
		if (main_genericstandalone_pcs_transmitpath_encoder_k) begin
			main_genericstandalone_pcs_transmitpath_encoder_alt7_rd0 <= 1'd1;
			main_genericstandalone_pcs_transmitpath_encoder_alt7_rd1 <= 1'd1;
		end
	end
	builder_a7_1000basex_transmitpath_state <= builder_a7_1000basex_transmitpath_next_state;
	if (main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value_ce) begin
		main_genericstandalone_pcs_transmitpath_c_type <= main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value;
	end
	main_genericstandalone_pcs_lp_abi_ping_o1 <= main_genericstandalone_pcs_lp_abi_ping_o0;
	if (main_genericstandalone_pcs_lp_abi_ping_o1) begin
		main_genericstandalone_pcs_lp_abi_o <= main_genericstandalone_pcs_lp_abi_obuffer;
	end
	main_genericstandalone_pcs_lp_abi_ping_toggle_o_r <= main_genericstandalone_pcs_lp_abi_ping_toggle_o;
	if (main_genericstandalone_pcs_lp_abi_pong_i) begin
		main_genericstandalone_pcs_lp_abi_pong_toggle_i <= (~main_genericstandalone_pcs_lp_abi_pong_toggle_i);
	end
	main_genericstandalone_pcs_seen_valid_ci_toggle_o_r <= main_genericstandalone_pcs_seen_valid_ci_toggle_o;
	main_genericstandalone_pcs_rx_config_reg_abi_toggle_o_r <= main_genericstandalone_pcs_rx_config_reg_abi_toggle_o;
	main_genericstandalone_pcs_rx_config_reg_ack_toggle_o_r <= main_genericstandalone_pcs_rx_config_reg_ack_toggle_o;
	if (main_genericstandalone_pcs_waittimer0_wait) begin
		if ((~main_genericstandalone_pcs_waittimer0_done)) begin
			main_genericstandalone_pcs_waittimer0_count <= (main_genericstandalone_pcs_waittimer0_count - 1'd1);
		end
	end else begin
		main_genericstandalone_pcs_waittimer0_count <= 21'd1250000;
	end
	if (main_genericstandalone_pcs_waittimer1_wait) begin
		if ((~main_genericstandalone_pcs_waittimer1_done)) begin
			main_genericstandalone_pcs_waittimer1_count <= (main_genericstandalone_pcs_waittimer1_count - 1'd1);
		end
	end else begin
		main_genericstandalone_pcs_waittimer1_count <= 18'd200000;
	end
	builder_a7_1000basex_fsm_state <= builder_a7_1000basex_fsm_next_state;
	if (main_genericstandalone_i) begin
		main_genericstandalone_toggle_i <= (~main_genericstandalone_toggle_i);
	end
	main_genericstandalone_buf <= {main_genericstandalone_tx_data1, main_genericstandalone_buf[19:10]};
	if (main_genericstandalone_tx_gap_inserter_counter_reset) begin
		main_genericstandalone_tx_gap_inserter_counter <= 1'd0;
	end else begin
		if (main_genericstandalone_tx_gap_inserter_counter_ce) begin
			main_genericstandalone_tx_gap_inserter_counter <= (main_genericstandalone_tx_gap_inserter_counter + 1'd1);
		end
	end
	builder_liteethmacgap_state <= builder_liteethmacgap_next_state;
	if (main_genericstandalone_preamble_inserter_clr_cnt) begin
		main_genericstandalone_preamble_inserter_cnt <= 1'd0;
	end else begin
		if (main_genericstandalone_preamble_inserter_inc_cnt) begin
			main_genericstandalone_preamble_inserter_cnt <= (main_genericstandalone_preamble_inserter_cnt + 1'd1);
		end
	end
	builder_liteethmacpreambleinserter_state <= builder_liteethmacpreambleinserter_next_state;
	if (main_genericstandalone_crc32_inserter_is_ongoing0) begin
		main_genericstandalone_crc32_inserter_cnt <= 2'd3;
	end else begin
		if ((main_genericstandalone_crc32_inserter_is_ongoing1 & (~main_genericstandalone_crc32_inserter_cnt_done))) begin
			main_genericstandalone_crc32_inserter_cnt <= (main_genericstandalone_crc32_inserter_cnt - main_genericstandalone_crc32_inserter_source_ack);
		end
	end
	if (main_genericstandalone_crc32_inserter_ce) begin
		main_genericstandalone_crc32_inserter_reg <= main_genericstandalone_crc32_inserter_next;
	end
	if (main_genericstandalone_crc32_inserter_reset) begin
		main_genericstandalone_crc32_inserter_reg <= 32'd4294967295;
	end
	builder_liteethmaccrc32inserter_state <= builder_liteethmaccrc32inserter_next_state;
	if (main_genericstandalone_padding_inserter_counter_reset) begin
		main_genericstandalone_padding_inserter_counter <= 1'd0;
	end else begin
		if (main_genericstandalone_padding_inserter_counter_ce) begin
			main_genericstandalone_padding_inserter_counter <= (main_genericstandalone_padding_inserter_counter + 1'd1);
		end
	end
	builder_liteethmacpaddinginserter_state <= builder_liteethmacpaddinginserter_next_state;
	if ((main_genericstandalone_tx_last_be_sink_stb & main_genericstandalone_tx_last_be_sink_ack)) begin
		if (main_genericstandalone_tx_last_be_sink_eop) begin
			main_genericstandalone_tx_last_be_ongoing <= 1'd1;
		end else begin
			if (main_genericstandalone_tx_last_be_sink_payload_last_be) begin
				main_genericstandalone_tx_last_be_ongoing <= 1'd0;
			end
		end
	end
	if ((main_genericstandalone_tx_converter_converter_source_stb & main_genericstandalone_tx_converter_converter_source_ack)) begin
		if (main_genericstandalone_tx_converter_converter_last) begin
			main_genericstandalone_tx_converter_converter_mux <= 1'd0;
		end else begin
			main_genericstandalone_tx_converter_converter_mux <= (main_genericstandalone_tx_converter_converter_mux + 1'd1);
		end
	end
	main_genericstandalone_tx_cdc_graycounter1_q_binary <= main_genericstandalone_tx_cdc_graycounter1_q_next_binary;
	main_genericstandalone_tx_cdc_graycounter1_q <= main_genericstandalone_tx_cdc_graycounter1_q_next;
	if (eth_tx_rst) begin
		main_genericstandalone_pcs_transmitpath_encoder2 <= 10'd0;
		main_genericstandalone_pcs_transmitpath_encoder3 <= 1'd0;
		main_genericstandalone_pcs_transmitpath_encoder_disp_in <= 1'd0;
		main_genericstandalone_pcs_transmitpath_encoder_code6b <= 6'd0;
		main_genericstandalone_pcs_transmitpath_encoder_code6b_unbalanced <= 1'd0;
		main_genericstandalone_pcs_transmitpath_encoder_code6b_flip <= 1'd0;
		main_genericstandalone_pcs_transmitpath_encoder_code4b <= 4'd0;
		main_genericstandalone_pcs_transmitpath_encoder_code4b_unbalanced <= 1'd0;
		main_genericstandalone_pcs_transmitpath_encoder_code4b_flip <= 1'd0;
		main_genericstandalone_pcs_transmitpath_encoder_alt7_rd0 <= 1'd0;
		main_genericstandalone_pcs_transmitpath_encoder_alt7_rd1 <= 1'd0;
		main_genericstandalone_pcs_transmitpath_parity <= 1'd0;
		main_genericstandalone_pcs_transmitpath_c_type <= 1'd0;
		main_genericstandalone_pcs_transmitpath_config_reg_buffer <= 16'd0;
		main_genericstandalone_pcs_transmitpath_timer <= 10'd0;
		main_genericstandalone_pcs_lp_abi_ping_o1 <= 1'd0;
		main_genericstandalone_pcs_checker_counter <= 20'd0;
		main_genericstandalone_pcs_checker_tick <= 1'd0;
		main_genericstandalone_pcs_checker_ok <= 1'd0;
		main_genericstandalone_pcs_waittimer0_count <= 21'd1250000;
		main_genericstandalone_pcs_waittimer1_count <= 18'd200000;
		main_genericstandalone_buf <= 20'd0;
		main_genericstandalone_tx_gap_inserter_counter <= 4'd0;
		main_genericstandalone_preamble_inserter_cnt <= 3'd0;
		main_genericstandalone_crc32_inserter_reg <= 32'd4294967295;
		main_genericstandalone_crc32_inserter_cnt <= 2'd3;
		main_genericstandalone_padding_inserter_counter <= 16'd1;
		main_genericstandalone_tx_last_be_ongoing <= 1'd1;
		main_genericstandalone_tx_converter_converter_mux <= 3'd0;
		main_genericstandalone_tx_cdc_graycounter1_q <= 7'd0;
		main_genericstandalone_tx_cdc_graycounter1_q_binary <= 7'd0;
		builder_a7_1000basex_transmitpath_state <= 3'd0;
		builder_a7_1000basex_fsm_state <= 3'd0;
		builder_liteethmacgap_state <= 1'd0;
		builder_liteethmacpreambleinserter_state <= 2'd0;
		builder_liteethmaccrc32inserter_state <= 2'd0;
		builder_liteethmacpaddinginserter_state <= 1'd0;
	end
	builder_xilinxmultiregimpl40 <= main_genericstandalone_pcs_lp_abi_ping_toggle_i;
	builder_xilinxmultiregimpl41 <= builder_xilinxmultiregimpl40;
	builder_xilinxmultiregimpl60 <= main_genericstandalone_pcs_lp_abi_ibuffer;
	builder_xilinxmultiregimpl61 <= builder_xilinxmultiregimpl60;
	builder_xilinxmultiregimpl70 <= main_genericstandalone_pcs_seen_valid_ci_toggle_i;
	builder_xilinxmultiregimpl71 <= builder_xilinxmultiregimpl70;
	builder_xilinxmultiregimpl80 <= main_genericstandalone_pcs_rx_config_reg_abi_toggle_i;
	builder_xilinxmultiregimpl81 <= builder_xilinxmultiregimpl80;
	builder_xilinxmultiregimpl90 <= main_genericstandalone_pcs_rx_config_reg_ack_toggle_i;
	builder_xilinxmultiregimpl91 <= builder_xilinxmultiregimpl90;
	builder_xilinxmultiregimpl150 <= main_genericstandalone_tx_cdc_graycounter0_q;
	builder_xilinxmultiregimpl151 <= builder_xilinxmultiregimpl150;
end

always @(posedge eth_tx_half_clk) begin
	main_genericstandalone_tx_data_half <= main_genericstandalone_buf;
end

always @(posedge icap_clk) begin
	main_genericstandalone_genericstandalone_icap_toggle_o_r <= main_genericstandalone_genericstandalone_icap_toggle_o;
	builder_icap_state <= builder_icap_next_state;
	if (main_genericstandalone_genericstandalone_icap_counter1_icap_next_value_ce) begin
		main_genericstandalone_genericstandalone_icap_counter1 <= main_genericstandalone_genericstandalone_icap_counter1_icap_next_value;
	end
	builder_xilinxmultiregimpl30 <= main_genericstandalone_genericstandalone_icap_toggle_i;
	builder_xilinxmultiregimpl31 <= builder_xilinxmultiregimpl30;
end

always @(posedge rio_clk) begin
	main_inout_8x0_inout_8x0_sample <= 1'd0;
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & main_inout_8x0_inout_8x0_ointerface0_address[1])) begin
		main_inout_8x0_inout_8x0_sensitivity <= main_inout_8x0_inout_8x0_ointerface0_data;
		if (main_inout_8x0_inout_8x0_ointerface0_address[0]) begin
			main_inout_8x0_inout_8x0_sample <= 1'd1;
		end
	end
	main_inout_8x1_inout_8x1_sample <= 1'd0;
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & main_inout_8x1_inout_8x1_ointerface1_address[1])) begin
		main_inout_8x1_inout_8x1_sensitivity <= main_inout_8x1_inout_8x1_ointerface1_data;
		if (main_inout_8x1_inout_8x1_ointerface1_address[0]) begin
			main_inout_8x1_inout_8x1_sample <= 1'd1;
		end
	end
	main_inout_8x2_inout_8x2_sample <= 1'd0;
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & main_inout_8x2_inout_8x2_ointerface2_address[1])) begin
		main_inout_8x2_inout_8x2_sensitivity <= main_inout_8x2_inout_8x2_ointerface2_data;
		if (main_inout_8x2_inout_8x2_ointerface2_address[0]) begin
			main_inout_8x2_inout_8x2_sample <= 1'd1;
		end
	end
	main_inout_8x3_inout_8x3_sample <= 1'd0;
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & main_inout_8x3_inout_8x3_ointerface3_address[1])) begin
		main_inout_8x3_inout_8x3_sensitivity <= main_inout_8x3_inout_8x3_ointerface3_data;
		if (main_inout_8x3_inout_8x3_ointerface3_address[0]) begin
			main_inout_8x3_inout_8x3_sample <= 1'd1;
		end
	end
	if (main_spimaster0_ointerface0_stb0) begin
		main_urukulmonitor0_current_address <= main_spimaster0_ointerface0_address0;
		main_urukulmonitor0_current_data <= main_spimaster0_ointerface0_data0;
		if ((main_spimaster0_ointerface0_address0 == 1'd1)) begin
			main_urukulmonitor0_cs <= main_spimaster0_ointerface0_data0[31:24];
			main_urukulmonitor0_data_length <= (main_spimaster0_ointerface0_data0[15:8] + 1'd1);
			main_urukulmonitor0_flags <= main_spimaster0_ointerface0_data0[7:0];
		end
	end
	if (main_spimaster1_ointerface1_stb0) begin
		main_urukulmonitor1_current_address <= main_spimaster1_ointerface1_address0;
		main_urukulmonitor1_current_data <= main_spimaster1_ointerface1_data0;
		if ((main_spimaster1_ointerface1_address0 == 1'd1)) begin
			main_urukulmonitor1_cs <= main_spimaster1_ointerface1_data0[31:24];
			main_urukulmonitor1_data_length <= (main_spimaster1_ointerface1_data0[15:8] + 1'd1);
			main_urukulmonitor1_flags <= main_spimaster1_ointerface1_data0[7:0];
		end
	end
	main_genericstandalone_rtio_core_sed_lane_dist_min_minus_timestamp <= (main_genericstandalone_rtio_core_sed_lane_dist_minimum_coarse_timestamp - main_genericstandalone_rtio_core_sed_lane_dist_coarse_timestamp);
	main_genericstandalone_rtio_core_sed_lane_dist_laneAmin_minus_timestamp <= (builder_sync_rhs_self3 - main_genericstandalone_rtio_core_sed_lane_dist_coarse_timestamp);
	main_genericstandalone_rtio_core_sed_lane_dist_laneBmin_minus_timestamp <= (builder_sync_rhs_self4 - main_genericstandalone_rtio_core_sed_lane_dist_coarse_timestamp);
	main_genericstandalone_rtio_core_sed_lane_dist_last_minus_timestamp <= (main_genericstandalone_rtio_core_sed_lane_dist_last_coarse_timestamp - main_genericstandalone_rtio_core_sed_lane_dist_coarse_timestamp);
	main_genericstandalone_rtio_core_sed_lane_dist_quash <= 1'd0;
	if ((main_genericstandalone_rtio_core_cri_chan_sel[15:0] == 6'd37)) begin
		main_genericstandalone_rtio_core_sed_lane_dist_quash <= 1'd1;
	end
	if (main_genericstandalone_rtio_core_sed_lane_dist_do_write) begin
		main_genericstandalone_rtio_core_sed_lane_dist_current_lane <= main_genericstandalone_rtio_core_sed_lane_dist_use_lanen;
		main_genericstandalone_rtio_core_sed_lane_dist_last_coarse_timestamp <= main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp[63:3];
		builder_sync_t_lhs_self = main_genericstandalone_rtio_core_sed_lane_dist_compensated_timestamp[63:3];
		case (main_genericstandalone_rtio_core_sed_lane_dist_use_lanen)
			1'd0: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps0 <= builder_sync_t_lhs_self;
			end
			1'd1: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps1 <= builder_sync_t_lhs_self;
			end
			2'd2: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps2 <= builder_sync_t_lhs_self;
			end
			2'd3: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps3 <= builder_sync_t_lhs_self;
			end
			3'd4: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps4 <= builder_sync_t_lhs_self;
			end
			3'd5: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps5 <= builder_sync_t_lhs_self;
			end
			3'd6: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps6 <= builder_sync_t_lhs_self;
			end
			3'd7: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps7 <= builder_sync_t_lhs_self;
			end
			4'd8: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps8 <= builder_sync_t_lhs_self;
			end
			4'd9: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps9 <= builder_sync_t_lhs_self;
			end
			4'd10: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps10 <= builder_sync_t_lhs_self;
			end
			4'd11: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps11 <= builder_sync_t_lhs_self;
			end
			4'd12: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps12 <= builder_sync_t_lhs_self;
			end
			4'd13: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps13 <= builder_sync_t_lhs_self;
			end
			4'd14: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps14 <= builder_sync_t_lhs_self;
			end
			default: begin
				main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps15 <= builder_sync_t_lhs_self;
			end
		endcase
		main_genericstandalone_rtio_core_sed_lane_dist_seqn <= (main_genericstandalone_rtio_core_sed_lane_dist_seqn + 1'd1);
	end
	if ((main_genericstandalone_rtio_core_cri_cmd == 1'd1)) begin
		main_genericstandalone_rtio_core_sed_lane_dist_o_status_underflow <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_sed_lane_dist_do_underflow) begin
		main_genericstandalone_rtio_core_sed_lane_dist_o_status_underflow <= 1'd1;
	end
	main_genericstandalone_rtio_core_sed_lane_dist_sequence_error <= main_genericstandalone_rtio_core_sed_lane_dist_do_sequence_error;
	main_genericstandalone_rtio_core_sed_lane_dist_sequence_error_channel <= main_genericstandalone_rtio_core_cri_chan_sel[15:0];
	if ((main_genericstandalone_rtio_core_sed_lane_dist_enable_spread & (main_genericstandalone_rtio_core_sed_lane_dist_current_lane_high_watermark | (~main_genericstandalone_rtio_core_sed_lane_dist_current_lane_writable)))) begin
		main_genericstandalone_rtio_core_sed_lane_dist_force_laneB <= 1'd1;
	end
	if (main_genericstandalone_rtio_core_sed_lane_dist_do_write) begin
		main_genericstandalone_rtio_core_sed_lane_dist_force_laneB <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered0_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered0_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_we & main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered0_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered0_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered0_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered0_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_we & main_genericstandalone_rtio_core_sed_syncfifobuffered0_syncfifo0_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered0_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered0_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered0_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered1_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered1_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_we & main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered1_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered1_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered1_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered1_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_we & main_genericstandalone_rtio_core_sed_syncfifobuffered1_syncfifo1_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered1_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered1_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered1_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered2_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered2_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_we & main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered2_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered2_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered2_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered2_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_we & main_genericstandalone_rtio_core_sed_syncfifobuffered2_syncfifo2_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered2_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered2_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered2_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered3_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered3_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_we & main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered3_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered3_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered3_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered3_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_we & main_genericstandalone_rtio_core_sed_syncfifobuffered3_syncfifo3_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered3_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered3_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered3_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered4_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered4_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_we & main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered4_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered4_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered4_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered4_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_we & main_genericstandalone_rtio_core_sed_syncfifobuffered4_syncfifo4_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered4_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered4_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered4_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered5_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered5_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_we & main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered5_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered5_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered5_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered5_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_we & main_genericstandalone_rtio_core_sed_syncfifobuffered5_syncfifo5_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered5_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered5_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered5_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered6_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered6_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_we & main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered6_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered6_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered6_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered6_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_we & main_genericstandalone_rtio_core_sed_syncfifobuffered6_syncfifo6_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered6_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered6_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered6_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered7_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered7_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_we & main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered7_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered7_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered7_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered7_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_we & main_genericstandalone_rtio_core_sed_syncfifobuffered7_syncfifo7_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered7_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered7_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered7_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered8_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered8_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_we & main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered8_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered8_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered8_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered8_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_we & main_genericstandalone_rtio_core_sed_syncfifobuffered8_syncfifo8_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered8_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered8_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered8_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered9_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered9_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_we & main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered9_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered9_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered9_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered9_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_we & main_genericstandalone_rtio_core_sed_syncfifobuffered9_syncfifo9_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered9_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered9_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered9_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered10_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered10_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_we & main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered10_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered10_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered10_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered10_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_we & main_genericstandalone_rtio_core_sed_syncfifobuffered10_syncfifo10_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered10_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered10_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered10_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered11_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered11_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_we & main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered11_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered11_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered11_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered11_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_we & main_genericstandalone_rtio_core_sed_syncfifobuffered11_syncfifo11_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered11_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered11_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered11_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered12_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered12_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_we & main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered12_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered12_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered12_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered12_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_we & main_genericstandalone_rtio_core_sed_syncfifobuffered12_syncfifo12_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered12_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered12_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered12_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered13_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered13_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_we & main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered13_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered13_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered13_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered13_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_we & main_genericstandalone_rtio_core_sed_syncfifobuffered13_syncfifo13_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered13_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered13_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered13_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered14_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered14_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_we & main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered14_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered14_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered14_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered14_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_we & main_genericstandalone_rtio_core_sed_syncfifobuffered14_syncfifo14_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered14_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered14_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered14_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_re) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered15_re) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered15_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_we & main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered15_replace))) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_produce <= (main_genericstandalone_rtio_core_sed_syncfifobuffered15_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered15_do_read) begin
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_consume <= (main_genericstandalone_rtio_core_sed_syncfifobuffered15_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_we & main_genericstandalone_rtio_core_sed_syncfifobuffered15_syncfifo15_writable) & (~main_genericstandalone_rtio_core_sed_syncfifobuffered15_replace))) begin
		if ((~main_genericstandalone_rtio_core_sed_syncfifobuffered15_do_read)) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_sed_syncfifobuffered15_do_read) begin
			main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 <= (main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 - 1'd1);
		end
	end
	main_genericstandalone_rtio_core_sed_gates_record16_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record0_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record16_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record0_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record16_payload_address <= main_genericstandalone_rtio_core_sed_gates_record0_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record16_payload_data <= main_genericstandalone_rtio_core_sed_gates_record0_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record16_seqn <= main_genericstandalone_rtio_core_sed_gates_record0_seqn;
	main_genericstandalone_rtio_core_sed_gates_record16_valid <= (main_genericstandalone_rtio_core_sed_gates_record0_re & main_genericstandalone_rtio_core_sed_gates_record0_readable);
	main_genericstandalone_rtio_core_sed_gates_record17_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record1_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record17_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record1_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record17_payload_address <= main_genericstandalone_rtio_core_sed_gates_record1_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record17_payload_data <= main_genericstandalone_rtio_core_sed_gates_record1_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record17_seqn <= main_genericstandalone_rtio_core_sed_gates_record1_seqn;
	main_genericstandalone_rtio_core_sed_gates_record17_valid <= (main_genericstandalone_rtio_core_sed_gates_record1_re & main_genericstandalone_rtio_core_sed_gates_record1_readable);
	main_genericstandalone_rtio_core_sed_gates_record18_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record2_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record18_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record2_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record18_payload_address <= main_genericstandalone_rtio_core_sed_gates_record2_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record18_payload_data <= main_genericstandalone_rtio_core_sed_gates_record2_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record18_seqn <= main_genericstandalone_rtio_core_sed_gates_record2_seqn;
	main_genericstandalone_rtio_core_sed_gates_record18_valid <= (main_genericstandalone_rtio_core_sed_gates_record2_re & main_genericstandalone_rtio_core_sed_gates_record2_readable);
	main_genericstandalone_rtio_core_sed_gates_record19_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record3_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record19_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record3_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record19_payload_address <= main_genericstandalone_rtio_core_sed_gates_record3_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record19_payload_data <= main_genericstandalone_rtio_core_sed_gates_record3_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record19_seqn <= main_genericstandalone_rtio_core_sed_gates_record3_seqn;
	main_genericstandalone_rtio_core_sed_gates_record19_valid <= (main_genericstandalone_rtio_core_sed_gates_record3_re & main_genericstandalone_rtio_core_sed_gates_record3_readable);
	main_genericstandalone_rtio_core_sed_gates_record20_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record4_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record20_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record4_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record20_payload_address <= main_genericstandalone_rtio_core_sed_gates_record4_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record20_payload_data <= main_genericstandalone_rtio_core_sed_gates_record4_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record20_seqn <= main_genericstandalone_rtio_core_sed_gates_record4_seqn;
	main_genericstandalone_rtio_core_sed_gates_record20_valid <= (main_genericstandalone_rtio_core_sed_gates_record4_re & main_genericstandalone_rtio_core_sed_gates_record4_readable);
	main_genericstandalone_rtio_core_sed_gates_record21_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record5_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record21_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record5_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record21_payload_address <= main_genericstandalone_rtio_core_sed_gates_record5_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record21_payload_data <= main_genericstandalone_rtio_core_sed_gates_record5_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record21_seqn <= main_genericstandalone_rtio_core_sed_gates_record5_seqn;
	main_genericstandalone_rtio_core_sed_gates_record21_valid <= (main_genericstandalone_rtio_core_sed_gates_record5_re & main_genericstandalone_rtio_core_sed_gates_record5_readable);
	main_genericstandalone_rtio_core_sed_gates_record22_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record6_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record22_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record6_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record22_payload_address <= main_genericstandalone_rtio_core_sed_gates_record6_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record22_payload_data <= main_genericstandalone_rtio_core_sed_gates_record6_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record22_seqn <= main_genericstandalone_rtio_core_sed_gates_record6_seqn;
	main_genericstandalone_rtio_core_sed_gates_record22_valid <= (main_genericstandalone_rtio_core_sed_gates_record6_re & main_genericstandalone_rtio_core_sed_gates_record6_readable);
	main_genericstandalone_rtio_core_sed_gates_record23_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record7_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record23_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record7_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record23_payload_address <= main_genericstandalone_rtio_core_sed_gates_record7_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record23_payload_data <= main_genericstandalone_rtio_core_sed_gates_record7_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record23_seqn <= main_genericstandalone_rtio_core_sed_gates_record7_seqn;
	main_genericstandalone_rtio_core_sed_gates_record23_valid <= (main_genericstandalone_rtio_core_sed_gates_record7_re & main_genericstandalone_rtio_core_sed_gates_record7_readable);
	main_genericstandalone_rtio_core_sed_gates_record24_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record8_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record24_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record8_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record24_payload_address <= main_genericstandalone_rtio_core_sed_gates_record8_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record24_payload_data <= main_genericstandalone_rtio_core_sed_gates_record8_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record24_seqn <= main_genericstandalone_rtio_core_sed_gates_record8_seqn;
	main_genericstandalone_rtio_core_sed_gates_record24_valid <= (main_genericstandalone_rtio_core_sed_gates_record8_re & main_genericstandalone_rtio_core_sed_gates_record8_readable);
	main_genericstandalone_rtio_core_sed_gates_record25_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record9_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record25_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record9_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record25_payload_address <= main_genericstandalone_rtio_core_sed_gates_record9_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record25_payload_data <= main_genericstandalone_rtio_core_sed_gates_record9_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record25_seqn <= main_genericstandalone_rtio_core_sed_gates_record9_seqn;
	main_genericstandalone_rtio_core_sed_gates_record25_valid <= (main_genericstandalone_rtio_core_sed_gates_record9_re & main_genericstandalone_rtio_core_sed_gates_record9_readable);
	main_genericstandalone_rtio_core_sed_gates_record26_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record10_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record26_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record10_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record26_payload_address <= main_genericstandalone_rtio_core_sed_gates_record10_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record26_payload_data <= main_genericstandalone_rtio_core_sed_gates_record10_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record26_seqn <= main_genericstandalone_rtio_core_sed_gates_record10_seqn;
	main_genericstandalone_rtio_core_sed_gates_record26_valid <= (main_genericstandalone_rtio_core_sed_gates_record10_re & main_genericstandalone_rtio_core_sed_gates_record10_readable);
	main_genericstandalone_rtio_core_sed_gates_record27_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record11_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record27_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record11_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record27_payload_address <= main_genericstandalone_rtio_core_sed_gates_record11_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record27_payload_data <= main_genericstandalone_rtio_core_sed_gates_record11_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record27_seqn <= main_genericstandalone_rtio_core_sed_gates_record11_seqn;
	main_genericstandalone_rtio_core_sed_gates_record27_valid <= (main_genericstandalone_rtio_core_sed_gates_record11_re & main_genericstandalone_rtio_core_sed_gates_record11_readable);
	main_genericstandalone_rtio_core_sed_gates_record28_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record12_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record28_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record12_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record28_payload_address <= main_genericstandalone_rtio_core_sed_gates_record12_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record28_payload_data <= main_genericstandalone_rtio_core_sed_gates_record12_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record28_seqn <= main_genericstandalone_rtio_core_sed_gates_record12_seqn;
	main_genericstandalone_rtio_core_sed_gates_record28_valid <= (main_genericstandalone_rtio_core_sed_gates_record12_re & main_genericstandalone_rtio_core_sed_gates_record12_readable);
	main_genericstandalone_rtio_core_sed_gates_record29_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record13_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record29_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record13_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record29_payload_address <= main_genericstandalone_rtio_core_sed_gates_record13_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record29_payload_data <= main_genericstandalone_rtio_core_sed_gates_record13_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record29_seqn <= main_genericstandalone_rtio_core_sed_gates_record13_seqn;
	main_genericstandalone_rtio_core_sed_gates_record29_valid <= (main_genericstandalone_rtio_core_sed_gates_record13_re & main_genericstandalone_rtio_core_sed_gates_record13_readable);
	main_genericstandalone_rtio_core_sed_gates_record30_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record14_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record30_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record14_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record30_payload_address <= main_genericstandalone_rtio_core_sed_gates_record14_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record30_payload_data <= main_genericstandalone_rtio_core_sed_gates_record14_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record30_seqn <= main_genericstandalone_rtio_core_sed_gates_record14_seqn;
	main_genericstandalone_rtio_core_sed_gates_record30_valid <= (main_genericstandalone_rtio_core_sed_gates_record14_re & main_genericstandalone_rtio_core_sed_gates_record14_readable);
	main_genericstandalone_rtio_core_sed_gates_record31_payload_channel <= main_genericstandalone_rtio_core_sed_gates_record15_payload_channel;
	main_genericstandalone_rtio_core_sed_gates_record31_payload_fine_ts <= main_genericstandalone_rtio_core_sed_gates_record15_payload_timestamp[2:0];
	main_genericstandalone_rtio_core_sed_gates_record31_payload_address <= main_genericstandalone_rtio_core_sed_gates_record15_payload_address;
	main_genericstandalone_rtio_core_sed_gates_record31_payload_data <= main_genericstandalone_rtio_core_sed_gates_record15_payload_data;
	main_genericstandalone_rtio_core_sed_gates_record31_seqn <= main_genericstandalone_rtio_core_sed_gates_record15_seqn;
	main_genericstandalone_rtio_core_sed_gates_record31_valid <= (main_genericstandalone_rtio_core_sed_gates_record15_re & main_genericstandalone_rtio_core_sed_gates_record15_readable);
	main_genericstandalone_rtio_core_sed_record0_valid1 <= main_genericstandalone_rtio_core_sed_record144_rec_valid;
	main_genericstandalone_rtio_core_sed_record0_payload_channel2 <= main_genericstandalone_rtio_core_sed_record144_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record144_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record0_payload_address2 <= main_genericstandalone_rtio_core_sed_record144_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record0_payload_data2 <= main_genericstandalone_rtio_core_sed_record144_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r0 <= main_genericstandalone_rtio_core_sed_record144_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r0 <= main_genericstandalone_rtio_core_sed_record144_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record1_valid1 <= main_genericstandalone_rtio_core_sed_record145_rec_valid;
	main_genericstandalone_rtio_core_sed_record1_payload_channel2 <= main_genericstandalone_rtio_core_sed_record145_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record145_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record1_payload_address2 <= main_genericstandalone_rtio_core_sed_record145_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record1_payload_data2 <= main_genericstandalone_rtio_core_sed_record145_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r1 <= main_genericstandalone_rtio_core_sed_record145_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r1 <= main_genericstandalone_rtio_core_sed_record145_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record2_valid1 <= main_genericstandalone_rtio_core_sed_record146_rec_valid;
	main_genericstandalone_rtio_core_sed_record2_payload_channel2 <= main_genericstandalone_rtio_core_sed_record146_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record146_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record2_payload_address2 <= main_genericstandalone_rtio_core_sed_record146_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record2_payload_data2 <= main_genericstandalone_rtio_core_sed_record146_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r2 <= main_genericstandalone_rtio_core_sed_record146_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r2 <= main_genericstandalone_rtio_core_sed_record146_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record3_valid1 <= main_genericstandalone_rtio_core_sed_record147_rec_valid;
	main_genericstandalone_rtio_core_sed_record3_payload_channel2 <= main_genericstandalone_rtio_core_sed_record147_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record147_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record3_payload_address2 <= main_genericstandalone_rtio_core_sed_record147_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record3_payload_data2 <= main_genericstandalone_rtio_core_sed_record147_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r3 <= main_genericstandalone_rtio_core_sed_record147_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r3 <= main_genericstandalone_rtio_core_sed_record147_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record4_valid1 <= main_genericstandalone_rtio_core_sed_record148_rec_valid;
	main_genericstandalone_rtio_core_sed_record4_payload_channel2 <= main_genericstandalone_rtio_core_sed_record148_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record148_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record4_payload_address2 <= main_genericstandalone_rtio_core_sed_record148_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record4_payload_data2 <= main_genericstandalone_rtio_core_sed_record148_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r4 <= main_genericstandalone_rtio_core_sed_record148_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r4 <= main_genericstandalone_rtio_core_sed_record148_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record5_valid1 <= main_genericstandalone_rtio_core_sed_record149_rec_valid;
	main_genericstandalone_rtio_core_sed_record5_payload_channel2 <= main_genericstandalone_rtio_core_sed_record149_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record149_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record5_payload_address2 <= main_genericstandalone_rtio_core_sed_record149_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record5_payload_data2 <= main_genericstandalone_rtio_core_sed_record149_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r5 <= main_genericstandalone_rtio_core_sed_record149_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r5 <= main_genericstandalone_rtio_core_sed_record149_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record6_valid1 <= main_genericstandalone_rtio_core_sed_record150_rec_valid;
	main_genericstandalone_rtio_core_sed_record6_payload_channel2 <= main_genericstandalone_rtio_core_sed_record150_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record150_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record6_payload_address2 <= main_genericstandalone_rtio_core_sed_record150_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record6_payload_data2 <= main_genericstandalone_rtio_core_sed_record150_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r6 <= main_genericstandalone_rtio_core_sed_record150_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r6 <= main_genericstandalone_rtio_core_sed_record150_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record7_valid1 <= main_genericstandalone_rtio_core_sed_record151_rec_valid;
	main_genericstandalone_rtio_core_sed_record7_payload_channel2 <= main_genericstandalone_rtio_core_sed_record151_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record151_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record7_payload_address2 <= main_genericstandalone_rtio_core_sed_record151_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record7_payload_data2 <= main_genericstandalone_rtio_core_sed_record151_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r7 <= main_genericstandalone_rtio_core_sed_record151_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r7 <= main_genericstandalone_rtio_core_sed_record151_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record8_valid1 <= main_genericstandalone_rtio_core_sed_record152_rec_valid;
	main_genericstandalone_rtio_core_sed_record8_payload_channel2 <= main_genericstandalone_rtio_core_sed_record152_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record152_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record8_payload_address2 <= main_genericstandalone_rtio_core_sed_record152_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record8_payload_data2 <= main_genericstandalone_rtio_core_sed_record152_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r8 <= main_genericstandalone_rtio_core_sed_record152_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r8 <= main_genericstandalone_rtio_core_sed_record152_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record9_valid1 <= main_genericstandalone_rtio_core_sed_record153_rec_valid;
	main_genericstandalone_rtio_core_sed_record9_payload_channel2 <= main_genericstandalone_rtio_core_sed_record153_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record153_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record9_payload_address2 <= main_genericstandalone_rtio_core_sed_record153_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record9_payload_data2 <= main_genericstandalone_rtio_core_sed_record153_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r9 <= main_genericstandalone_rtio_core_sed_record153_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r9 <= main_genericstandalone_rtio_core_sed_record153_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record10_valid1 <= main_genericstandalone_rtio_core_sed_record154_rec_valid;
	main_genericstandalone_rtio_core_sed_record10_payload_channel2 <= main_genericstandalone_rtio_core_sed_record154_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record154_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record10_payload_address2 <= main_genericstandalone_rtio_core_sed_record154_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record10_payload_data2 <= main_genericstandalone_rtio_core_sed_record154_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r10 <= main_genericstandalone_rtio_core_sed_record154_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r10 <= main_genericstandalone_rtio_core_sed_record154_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record11_valid1 <= main_genericstandalone_rtio_core_sed_record155_rec_valid;
	main_genericstandalone_rtio_core_sed_record11_payload_channel2 <= main_genericstandalone_rtio_core_sed_record155_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record155_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record11_payload_address2 <= main_genericstandalone_rtio_core_sed_record155_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record11_payload_data2 <= main_genericstandalone_rtio_core_sed_record155_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r11 <= main_genericstandalone_rtio_core_sed_record155_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r11 <= main_genericstandalone_rtio_core_sed_record155_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record12_valid1 <= main_genericstandalone_rtio_core_sed_record156_rec_valid;
	main_genericstandalone_rtio_core_sed_record12_payload_channel2 <= main_genericstandalone_rtio_core_sed_record156_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record156_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record12_payload_address2 <= main_genericstandalone_rtio_core_sed_record156_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record12_payload_data2 <= main_genericstandalone_rtio_core_sed_record156_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r12 <= main_genericstandalone_rtio_core_sed_record156_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r12 <= main_genericstandalone_rtio_core_sed_record156_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record13_valid1 <= main_genericstandalone_rtio_core_sed_record157_rec_valid;
	main_genericstandalone_rtio_core_sed_record13_payload_channel2 <= main_genericstandalone_rtio_core_sed_record157_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record157_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record13_payload_address2 <= main_genericstandalone_rtio_core_sed_record157_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record13_payload_data2 <= main_genericstandalone_rtio_core_sed_record157_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r13 <= main_genericstandalone_rtio_core_sed_record157_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r13 <= main_genericstandalone_rtio_core_sed_record157_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record14_valid1 <= main_genericstandalone_rtio_core_sed_record158_rec_valid;
	main_genericstandalone_rtio_core_sed_record14_payload_channel2 <= main_genericstandalone_rtio_core_sed_record158_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record158_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record14_payload_address2 <= main_genericstandalone_rtio_core_sed_record158_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record14_payload_data2 <= main_genericstandalone_rtio_core_sed_record158_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r14 <= main_genericstandalone_rtio_core_sed_record158_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r14 <= main_genericstandalone_rtio_core_sed_record158_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record15_valid1 <= main_genericstandalone_rtio_core_sed_record159_rec_valid;
	main_genericstandalone_rtio_core_sed_record15_payload_channel2 <= main_genericstandalone_rtio_core_sed_record159_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1 <= main_genericstandalone_rtio_core_sed_record159_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record15_payload_address2 <= main_genericstandalone_rtio_core_sed_record159_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record15_payload_data2 <= main_genericstandalone_rtio_core_sed_record159_rec_payload_data;
	main_genericstandalone_rtio_core_sed_replace_occured_r15 <= main_genericstandalone_rtio_core_sed_record159_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_nondata_replace_occured_r15 <= main_genericstandalone_rtio_core_sed_record159_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_collision <= 1'd0;
	main_genericstandalone_rtio_core_sed_collision_channel <= 1'd0;
	if ((main_genericstandalone_rtio_core_sed_record0_valid1 & main_genericstandalone_rtio_core_sed_record0_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record0_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record1_valid1 & main_genericstandalone_rtio_core_sed_record1_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record1_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record2_valid1 & main_genericstandalone_rtio_core_sed_record2_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record2_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record3_valid1 & main_genericstandalone_rtio_core_sed_record3_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record3_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record4_valid1 & main_genericstandalone_rtio_core_sed_record4_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record4_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record5_valid1 & main_genericstandalone_rtio_core_sed_record5_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record5_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record6_valid1 & main_genericstandalone_rtio_core_sed_record6_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record6_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record7_valid1 & main_genericstandalone_rtio_core_sed_record7_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record7_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record8_valid1 & main_genericstandalone_rtio_core_sed_record8_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record8_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record9_valid1 & main_genericstandalone_rtio_core_sed_record9_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record9_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record10_valid1 & main_genericstandalone_rtio_core_sed_record10_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record10_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record11_valid1 & main_genericstandalone_rtio_core_sed_record11_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record11_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record12_valid1 & main_genericstandalone_rtio_core_sed_record12_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record12_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record13_valid1 & main_genericstandalone_rtio_core_sed_record13_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record13_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record14_valid1 & main_genericstandalone_rtio_core_sed_record14_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record14_payload_channel2;
	end
	if ((main_genericstandalone_rtio_core_sed_record15_valid1 & main_genericstandalone_rtio_core_sed_record15_collision)) begin
		main_genericstandalone_rtio_core_sed_collision <= 1'd1;
		main_genericstandalone_rtio_core_sed_collision_channel <= main_genericstandalone_rtio_core_sed_record15_payload_channel2;
	end
	main_inout_8x0_inout_8x0_ointerface0_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected0 | main_genericstandalone_rtio_core_sed_selected1) | main_genericstandalone_rtio_core_sed_selected2) | main_genericstandalone_rtio_core_sed_selected3) | main_genericstandalone_rtio_core_sed_selected4) | main_genericstandalone_rtio_core_sed_selected5) | main_genericstandalone_rtio_core_sed_selected6) | main_genericstandalone_rtio_core_sed_selected7) | main_genericstandalone_rtio_core_sed_selected8) | main_genericstandalone_rtio_core_sed_selected9) | main_genericstandalone_rtio_core_sed_selected10) | main_genericstandalone_rtio_core_sed_selected11) | main_genericstandalone_rtio_core_sed_selected12) | main_genericstandalone_rtio_core_sed_selected13) | main_genericstandalone_rtio_core_sed_selected14) | main_genericstandalone_rtio_core_sed_selected15);
	main_inout_8x0_inout_8x0_ointerface0_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected0 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected1 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected2 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected3 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected4 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected5 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected6 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected7 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected8 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected9 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected10 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected11 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected12 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected13 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected14 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected15 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x0_inout_8x0_ointerface0_address <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected0 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected1 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected2 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected3 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected4 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected5 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected6 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected7 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected8 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected9 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected10 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected11 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected12 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected13 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected14 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected15 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_inout_8x0_inout_8x0_ointerface0_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected0 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected1 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected2 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected3 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected4 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected5 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected6 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected7 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected8 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected9 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected10 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected11 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected12 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected13 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected14 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected15 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected16 | main_genericstandalone_rtio_core_sed_selected17) | main_genericstandalone_rtio_core_sed_selected18) | main_genericstandalone_rtio_core_sed_selected19) | main_genericstandalone_rtio_core_sed_selected20) | main_genericstandalone_rtio_core_sed_selected21) | main_genericstandalone_rtio_core_sed_selected22) | main_genericstandalone_rtio_core_sed_selected23) | main_genericstandalone_rtio_core_sed_selected24) | main_genericstandalone_rtio_core_sed_selected25) | main_genericstandalone_rtio_core_sed_selected26) | main_genericstandalone_rtio_core_sed_selected27) | main_genericstandalone_rtio_core_sed_selected28) | main_genericstandalone_rtio_core_sed_selected29) | main_genericstandalone_rtio_core_sed_selected30) | main_genericstandalone_rtio_core_sed_selected31);
	main_inout_8x1_inout_8x1_ointerface1_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected16 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected17 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected18 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected19 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected20 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected21 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected22 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected23 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected24 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected25 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected26 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected27 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected28 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected29 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected30 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected31 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_address <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected16 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected17 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected18 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected19 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected20 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected21 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected22 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected23 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected24 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected25 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected26 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected27 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected28 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected29 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected30 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected31 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected16 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected17 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected18 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected19 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected20 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected21 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected22 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected23 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected24 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected25 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected26 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected27 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected28 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected29 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected30 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected31 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected32 | main_genericstandalone_rtio_core_sed_selected33) | main_genericstandalone_rtio_core_sed_selected34) | main_genericstandalone_rtio_core_sed_selected35) | main_genericstandalone_rtio_core_sed_selected36) | main_genericstandalone_rtio_core_sed_selected37) | main_genericstandalone_rtio_core_sed_selected38) | main_genericstandalone_rtio_core_sed_selected39) | main_genericstandalone_rtio_core_sed_selected40) | main_genericstandalone_rtio_core_sed_selected41) | main_genericstandalone_rtio_core_sed_selected42) | main_genericstandalone_rtio_core_sed_selected43) | main_genericstandalone_rtio_core_sed_selected44) | main_genericstandalone_rtio_core_sed_selected45) | main_genericstandalone_rtio_core_sed_selected46) | main_genericstandalone_rtio_core_sed_selected47);
	main_inout_8x2_inout_8x2_ointerface2_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected32 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected33 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected34 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected35 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected36 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected37 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected38 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected39 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected40 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected41 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected42 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected43 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected44 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected45 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected46 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected47 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_address <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected32 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected33 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected34 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected35 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected36 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected37 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected38 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected39 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected40 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected41 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected42 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected43 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected44 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected45 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected46 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected47 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected32 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected33 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected34 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected35 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected36 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected37 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected38 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected39 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected40 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected41 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected42 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected43 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected44 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected45 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected46 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected47 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected48 | main_genericstandalone_rtio_core_sed_selected49) | main_genericstandalone_rtio_core_sed_selected50) | main_genericstandalone_rtio_core_sed_selected51) | main_genericstandalone_rtio_core_sed_selected52) | main_genericstandalone_rtio_core_sed_selected53) | main_genericstandalone_rtio_core_sed_selected54) | main_genericstandalone_rtio_core_sed_selected55) | main_genericstandalone_rtio_core_sed_selected56) | main_genericstandalone_rtio_core_sed_selected57) | main_genericstandalone_rtio_core_sed_selected58) | main_genericstandalone_rtio_core_sed_selected59) | main_genericstandalone_rtio_core_sed_selected60) | main_genericstandalone_rtio_core_sed_selected61) | main_genericstandalone_rtio_core_sed_selected62) | main_genericstandalone_rtio_core_sed_selected63);
	main_inout_8x3_inout_8x3_ointerface3_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected48 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected49 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected50 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected51 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected52 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected53 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected54 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected55 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected56 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected57 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected58 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected59 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected60 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected61 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected62 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected63 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_address <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected48 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected49 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected50 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected51 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected52 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected53 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected54 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected55 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected56 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected57 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected58 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected59 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected60 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected61 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected62 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected63 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected48 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected49 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected50 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected51 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected52 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected53 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected54 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected55 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected56 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected57 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected58 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected59 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected60 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected61 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected62 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected63 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x0_stb0 <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected64 | main_genericstandalone_rtio_core_sed_selected65) | main_genericstandalone_rtio_core_sed_selected66) | main_genericstandalone_rtio_core_sed_selected67) | main_genericstandalone_rtio_core_sed_selected68) | main_genericstandalone_rtio_core_sed_selected69) | main_genericstandalone_rtio_core_sed_selected70) | main_genericstandalone_rtio_core_sed_selected71) | main_genericstandalone_rtio_core_sed_selected72) | main_genericstandalone_rtio_core_sed_selected73) | main_genericstandalone_rtio_core_sed_selected74) | main_genericstandalone_rtio_core_sed_selected75) | main_genericstandalone_rtio_core_sed_selected76) | main_genericstandalone_rtio_core_sed_selected77) | main_genericstandalone_rtio_core_sed_selected78) | main_genericstandalone_rtio_core_sed_selected79);
	main_output_8x0_fine_ts0 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected64 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected65 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected66 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected67 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected68 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected69 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected70 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected71 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected72 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected73 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected74 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected75 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected76 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected77 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected78 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected79 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x0_data0 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected64 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected65 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected66 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected67 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected68 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected69 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected70 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected71 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected72 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected73 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected74 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected75 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected76 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected77 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected78 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected79 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x1_stb0 <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected80 | main_genericstandalone_rtio_core_sed_selected81) | main_genericstandalone_rtio_core_sed_selected82) | main_genericstandalone_rtio_core_sed_selected83) | main_genericstandalone_rtio_core_sed_selected84) | main_genericstandalone_rtio_core_sed_selected85) | main_genericstandalone_rtio_core_sed_selected86) | main_genericstandalone_rtio_core_sed_selected87) | main_genericstandalone_rtio_core_sed_selected88) | main_genericstandalone_rtio_core_sed_selected89) | main_genericstandalone_rtio_core_sed_selected90) | main_genericstandalone_rtio_core_sed_selected91) | main_genericstandalone_rtio_core_sed_selected92) | main_genericstandalone_rtio_core_sed_selected93) | main_genericstandalone_rtio_core_sed_selected94) | main_genericstandalone_rtio_core_sed_selected95);
	main_output_8x1_fine_ts0 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected80 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected81 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected82 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected83 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected84 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected85 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected86 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected87 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected88 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected89 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected90 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected91 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected92 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected93 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected94 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected95 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x1_data0 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected80 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected81 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected82 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected83 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected84 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected85 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected86 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected87 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected88 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected89 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected90 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected91 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected92 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected93 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected94 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected95 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x2_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected96 | main_genericstandalone_rtio_core_sed_selected97) | main_genericstandalone_rtio_core_sed_selected98) | main_genericstandalone_rtio_core_sed_selected99) | main_genericstandalone_rtio_core_sed_selected100) | main_genericstandalone_rtio_core_sed_selected101) | main_genericstandalone_rtio_core_sed_selected102) | main_genericstandalone_rtio_core_sed_selected103) | main_genericstandalone_rtio_core_sed_selected104) | main_genericstandalone_rtio_core_sed_selected105) | main_genericstandalone_rtio_core_sed_selected106) | main_genericstandalone_rtio_core_sed_selected107) | main_genericstandalone_rtio_core_sed_selected108) | main_genericstandalone_rtio_core_sed_selected109) | main_genericstandalone_rtio_core_sed_selected110) | main_genericstandalone_rtio_core_sed_selected111);
	main_output_8x2_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected96 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected97 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected98 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected99 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected100 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected101 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected102 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected103 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected104 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected105 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected106 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected107 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected108 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected109 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected110 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected111 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x2_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected96 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected97 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected98 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected99 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected100 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected101 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected102 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected103 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected104 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected105 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected106 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected107 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected108 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected109 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected110 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected111 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x3_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected112 | main_genericstandalone_rtio_core_sed_selected113) | main_genericstandalone_rtio_core_sed_selected114) | main_genericstandalone_rtio_core_sed_selected115) | main_genericstandalone_rtio_core_sed_selected116) | main_genericstandalone_rtio_core_sed_selected117) | main_genericstandalone_rtio_core_sed_selected118) | main_genericstandalone_rtio_core_sed_selected119) | main_genericstandalone_rtio_core_sed_selected120) | main_genericstandalone_rtio_core_sed_selected121) | main_genericstandalone_rtio_core_sed_selected122) | main_genericstandalone_rtio_core_sed_selected123) | main_genericstandalone_rtio_core_sed_selected124) | main_genericstandalone_rtio_core_sed_selected125) | main_genericstandalone_rtio_core_sed_selected126) | main_genericstandalone_rtio_core_sed_selected127);
	main_output_8x3_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected112 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected113 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected114 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected115 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected116 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected117 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected118 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected119 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected120 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected121 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected122 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected123 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected124 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected125 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected126 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected127 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x3_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected112 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected113 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected114 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected115 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected116 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected117 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected118 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected119 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected120 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected121 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected122 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected123 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected124 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected125 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected126 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected127 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x4_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected128 | main_genericstandalone_rtio_core_sed_selected129) | main_genericstandalone_rtio_core_sed_selected130) | main_genericstandalone_rtio_core_sed_selected131) | main_genericstandalone_rtio_core_sed_selected132) | main_genericstandalone_rtio_core_sed_selected133) | main_genericstandalone_rtio_core_sed_selected134) | main_genericstandalone_rtio_core_sed_selected135) | main_genericstandalone_rtio_core_sed_selected136) | main_genericstandalone_rtio_core_sed_selected137) | main_genericstandalone_rtio_core_sed_selected138) | main_genericstandalone_rtio_core_sed_selected139) | main_genericstandalone_rtio_core_sed_selected140) | main_genericstandalone_rtio_core_sed_selected141) | main_genericstandalone_rtio_core_sed_selected142) | main_genericstandalone_rtio_core_sed_selected143);
	main_output_8x4_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected128 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected129 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected130 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected131 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected132 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected133 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected134 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected135 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected136 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected137 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected138 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected139 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected140 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected141 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected142 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected143 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x4_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected128 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected129 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected130 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected131 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected132 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected133 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected134 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected135 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected136 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected137 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected138 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected139 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected140 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected141 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected142 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected143 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x5_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected144 | main_genericstandalone_rtio_core_sed_selected145) | main_genericstandalone_rtio_core_sed_selected146) | main_genericstandalone_rtio_core_sed_selected147) | main_genericstandalone_rtio_core_sed_selected148) | main_genericstandalone_rtio_core_sed_selected149) | main_genericstandalone_rtio_core_sed_selected150) | main_genericstandalone_rtio_core_sed_selected151) | main_genericstandalone_rtio_core_sed_selected152) | main_genericstandalone_rtio_core_sed_selected153) | main_genericstandalone_rtio_core_sed_selected154) | main_genericstandalone_rtio_core_sed_selected155) | main_genericstandalone_rtio_core_sed_selected156) | main_genericstandalone_rtio_core_sed_selected157) | main_genericstandalone_rtio_core_sed_selected158) | main_genericstandalone_rtio_core_sed_selected159);
	main_output_8x5_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected144 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected145 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected146 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected147 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected148 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected149 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected150 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected151 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected152 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected153 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected154 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected155 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected156 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected157 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected158 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected159 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x5_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected144 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected145 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected146 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected147 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected148 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected149 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected150 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected151 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected152 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected153 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected154 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected155 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected156 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected157 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected158 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected159 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x6_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected160 | main_genericstandalone_rtio_core_sed_selected161) | main_genericstandalone_rtio_core_sed_selected162) | main_genericstandalone_rtio_core_sed_selected163) | main_genericstandalone_rtio_core_sed_selected164) | main_genericstandalone_rtio_core_sed_selected165) | main_genericstandalone_rtio_core_sed_selected166) | main_genericstandalone_rtio_core_sed_selected167) | main_genericstandalone_rtio_core_sed_selected168) | main_genericstandalone_rtio_core_sed_selected169) | main_genericstandalone_rtio_core_sed_selected170) | main_genericstandalone_rtio_core_sed_selected171) | main_genericstandalone_rtio_core_sed_selected172) | main_genericstandalone_rtio_core_sed_selected173) | main_genericstandalone_rtio_core_sed_selected174) | main_genericstandalone_rtio_core_sed_selected175);
	main_output_8x6_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected160 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected161 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected162 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected163 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected164 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected165 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected166 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected167 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected168 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected169 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected170 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected171 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected172 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected173 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected174 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected175 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x6_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected160 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected161 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected162 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected163 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected164 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected165 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected166 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected167 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected168 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected169 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected170 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected171 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected172 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected173 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected174 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected175 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x7_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected176 | main_genericstandalone_rtio_core_sed_selected177) | main_genericstandalone_rtio_core_sed_selected178) | main_genericstandalone_rtio_core_sed_selected179) | main_genericstandalone_rtio_core_sed_selected180) | main_genericstandalone_rtio_core_sed_selected181) | main_genericstandalone_rtio_core_sed_selected182) | main_genericstandalone_rtio_core_sed_selected183) | main_genericstandalone_rtio_core_sed_selected184) | main_genericstandalone_rtio_core_sed_selected185) | main_genericstandalone_rtio_core_sed_selected186) | main_genericstandalone_rtio_core_sed_selected187) | main_genericstandalone_rtio_core_sed_selected188) | main_genericstandalone_rtio_core_sed_selected189) | main_genericstandalone_rtio_core_sed_selected190) | main_genericstandalone_rtio_core_sed_selected191);
	main_output_8x7_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected176 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected177 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected178 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected179 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected180 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected181 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected182 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected183 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected184 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected185 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected186 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected187 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected188 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected189 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected190 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected191 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x7_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected176 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected177 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected178 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected179 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected180 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected181 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected182 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected183 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected184 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected185 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected186 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected187 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected188 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected189 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected190 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected191 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x8_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected192 | main_genericstandalone_rtio_core_sed_selected193) | main_genericstandalone_rtio_core_sed_selected194) | main_genericstandalone_rtio_core_sed_selected195) | main_genericstandalone_rtio_core_sed_selected196) | main_genericstandalone_rtio_core_sed_selected197) | main_genericstandalone_rtio_core_sed_selected198) | main_genericstandalone_rtio_core_sed_selected199) | main_genericstandalone_rtio_core_sed_selected200) | main_genericstandalone_rtio_core_sed_selected201) | main_genericstandalone_rtio_core_sed_selected202) | main_genericstandalone_rtio_core_sed_selected203) | main_genericstandalone_rtio_core_sed_selected204) | main_genericstandalone_rtio_core_sed_selected205) | main_genericstandalone_rtio_core_sed_selected206) | main_genericstandalone_rtio_core_sed_selected207);
	main_output_8x8_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected192 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected193 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected194 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected195 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected196 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected197 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected198 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected199 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected200 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected201 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected202 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected203 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected204 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected205 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected206 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected207 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x8_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected192 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected193 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected194 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected195 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected196 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected197 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected198 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected199 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected200 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected201 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected202 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected203 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected204 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected205 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected206 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected207 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x9_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected208 | main_genericstandalone_rtio_core_sed_selected209) | main_genericstandalone_rtio_core_sed_selected210) | main_genericstandalone_rtio_core_sed_selected211) | main_genericstandalone_rtio_core_sed_selected212) | main_genericstandalone_rtio_core_sed_selected213) | main_genericstandalone_rtio_core_sed_selected214) | main_genericstandalone_rtio_core_sed_selected215) | main_genericstandalone_rtio_core_sed_selected216) | main_genericstandalone_rtio_core_sed_selected217) | main_genericstandalone_rtio_core_sed_selected218) | main_genericstandalone_rtio_core_sed_selected219) | main_genericstandalone_rtio_core_sed_selected220) | main_genericstandalone_rtio_core_sed_selected221) | main_genericstandalone_rtio_core_sed_selected222) | main_genericstandalone_rtio_core_sed_selected223);
	main_output_8x9_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected208 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected209 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected210 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected211 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected212 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected213 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected214 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected215 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected216 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected217 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected218 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected219 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected220 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected221 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected222 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected223 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x9_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected208 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected209 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected210 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected211 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected212 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected213 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected214 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected215 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected216 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected217 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected218 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected219 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected220 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected221 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected222 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected223 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x10_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected224 | main_genericstandalone_rtio_core_sed_selected225) | main_genericstandalone_rtio_core_sed_selected226) | main_genericstandalone_rtio_core_sed_selected227) | main_genericstandalone_rtio_core_sed_selected228) | main_genericstandalone_rtio_core_sed_selected229) | main_genericstandalone_rtio_core_sed_selected230) | main_genericstandalone_rtio_core_sed_selected231) | main_genericstandalone_rtio_core_sed_selected232) | main_genericstandalone_rtio_core_sed_selected233) | main_genericstandalone_rtio_core_sed_selected234) | main_genericstandalone_rtio_core_sed_selected235) | main_genericstandalone_rtio_core_sed_selected236) | main_genericstandalone_rtio_core_sed_selected237) | main_genericstandalone_rtio_core_sed_selected238) | main_genericstandalone_rtio_core_sed_selected239);
	main_output_8x10_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected224 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected225 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected226 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected227 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected228 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected229 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected230 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected231 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected232 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected233 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected234 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected235 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected236 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected237 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected238 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected239 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x10_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected224 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected225 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected226 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected227 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected228 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected229 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected230 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected231 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected232 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected233 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected234 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected235 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected236 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected237 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected238 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected239 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x11_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected240 | main_genericstandalone_rtio_core_sed_selected241) | main_genericstandalone_rtio_core_sed_selected242) | main_genericstandalone_rtio_core_sed_selected243) | main_genericstandalone_rtio_core_sed_selected244) | main_genericstandalone_rtio_core_sed_selected245) | main_genericstandalone_rtio_core_sed_selected246) | main_genericstandalone_rtio_core_sed_selected247) | main_genericstandalone_rtio_core_sed_selected248) | main_genericstandalone_rtio_core_sed_selected249) | main_genericstandalone_rtio_core_sed_selected250) | main_genericstandalone_rtio_core_sed_selected251) | main_genericstandalone_rtio_core_sed_selected252) | main_genericstandalone_rtio_core_sed_selected253) | main_genericstandalone_rtio_core_sed_selected254) | main_genericstandalone_rtio_core_sed_selected255);
	main_output_8x11_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected240 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected241 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected242 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected243 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected244 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected245 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected246 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected247 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected248 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected249 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected250 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected251 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected252 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected253 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected254 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected255 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x11_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected240 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected241 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected242 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected243 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected244 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected245 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected246 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected247 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected248 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected249 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected250 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected251 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected252 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected253 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected254 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected255 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_spimaster0_ointerface0_stb0 <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected256 | main_genericstandalone_rtio_core_sed_selected257) | main_genericstandalone_rtio_core_sed_selected258) | main_genericstandalone_rtio_core_sed_selected259) | main_genericstandalone_rtio_core_sed_selected260) | main_genericstandalone_rtio_core_sed_selected261) | main_genericstandalone_rtio_core_sed_selected262) | main_genericstandalone_rtio_core_sed_selected263) | main_genericstandalone_rtio_core_sed_selected264) | main_genericstandalone_rtio_core_sed_selected265) | main_genericstandalone_rtio_core_sed_selected266) | main_genericstandalone_rtio_core_sed_selected267) | main_genericstandalone_rtio_core_sed_selected268) | main_genericstandalone_rtio_core_sed_selected269) | main_genericstandalone_rtio_core_sed_selected270) | main_genericstandalone_rtio_core_sed_selected271);
	main_spimaster0_ointerface0_address0 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected256 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected257 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected258 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected259 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected260 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected261 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected262 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected263 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected264 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected265 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected266 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected267 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected268 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected269 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected270 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected271 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_spimaster0_ointerface0_data0 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected256 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected257 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected258 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected259 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected260 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected261 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected262 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected263 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected264 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected265 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected266 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected267 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected268 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected269 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected270 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected271 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x0_stb1 <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected272 | main_genericstandalone_rtio_core_sed_selected273) | main_genericstandalone_rtio_core_sed_selected274) | main_genericstandalone_rtio_core_sed_selected275) | main_genericstandalone_rtio_core_sed_selected276) | main_genericstandalone_rtio_core_sed_selected277) | main_genericstandalone_rtio_core_sed_selected278) | main_genericstandalone_rtio_core_sed_selected279) | main_genericstandalone_rtio_core_sed_selected280) | main_genericstandalone_rtio_core_sed_selected281) | main_genericstandalone_rtio_core_sed_selected282) | main_genericstandalone_rtio_core_sed_selected283) | main_genericstandalone_rtio_core_sed_selected284) | main_genericstandalone_rtio_core_sed_selected285) | main_genericstandalone_rtio_core_sed_selected286) | main_genericstandalone_rtio_core_sed_selected287);
	main_output_8x0_fine_ts1 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected272 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected273 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected274 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected275 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected276 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected277 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected278 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected279 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected280 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected281 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected282 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected283 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected284 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected285 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected286 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected287 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x0_data1 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected272 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected273 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected274 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected275 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected276 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected277 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected278 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected279 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected280 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected281 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected282 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected283 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected284 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected285 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected286 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected287 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x12_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected288 | main_genericstandalone_rtio_core_sed_selected289) | main_genericstandalone_rtio_core_sed_selected290) | main_genericstandalone_rtio_core_sed_selected291) | main_genericstandalone_rtio_core_sed_selected292) | main_genericstandalone_rtio_core_sed_selected293) | main_genericstandalone_rtio_core_sed_selected294) | main_genericstandalone_rtio_core_sed_selected295) | main_genericstandalone_rtio_core_sed_selected296) | main_genericstandalone_rtio_core_sed_selected297) | main_genericstandalone_rtio_core_sed_selected298) | main_genericstandalone_rtio_core_sed_selected299) | main_genericstandalone_rtio_core_sed_selected300) | main_genericstandalone_rtio_core_sed_selected301) | main_genericstandalone_rtio_core_sed_selected302) | main_genericstandalone_rtio_core_sed_selected303);
	main_output_8x12_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected288 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected289 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected290 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected291 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected292 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected293 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected294 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected295 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected296 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected297 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected298 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected299 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected300 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected301 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected302 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected303 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x12_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected288 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected289 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected290 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected291 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected292 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected293 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected294 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected295 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected296 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected297 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected298 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected299 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected300 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected301 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected302 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected303 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x13_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected304 | main_genericstandalone_rtio_core_sed_selected305) | main_genericstandalone_rtio_core_sed_selected306) | main_genericstandalone_rtio_core_sed_selected307) | main_genericstandalone_rtio_core_sed_selected308) | main_genericstandalone_rtio_core_sed_selected309) | main_genericstandalone_rtio_core_sed_selected310) | main_genericstandalone_rtio_core_sed_selected311) | main_genericstandalone_rtio_core_sed_selected312) | main_genericstandalone_rtio_core_sed_selected313) | main_genericstandalone_rtio_core_sed_selected314) | main_genericstandalone_rtio_core_sed_selected315) | main_genericstandalone_rtio_core_sed_selected316) | main_genericstandalone_rtio_core_sed_selected317) | main_genericstandalone_rtio_core_sed_selected318) | main_genericstandalone_rtio_core_sed_selected319);
	main_output_8x13_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected304 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected305 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected306 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected307 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected308 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected309 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected310 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected311 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected312 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected313 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected314 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected315 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected316 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected317 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected318 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected319 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x13_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected304 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected305 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected306 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected307 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected308 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected309 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected310 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected311 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected312 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected313 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected314 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected315 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected316 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected317 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected318 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected319 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x14_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected320 | main_genericstandalone_rtio_core_sed_selected321) | main_genericstandalone_rtio_core_sed_selected322) | main_genericstandalone_rtio_core_sed_selected323) | main_genericstandalone_rtio_core_sed_selected324) | main_genericstandalone_rtio_core_sed_selected325) | main_genericstandalone_rtio_core_sed_selected326) | main_genericstandalone_rtio_core_sed_selected327) | main_genericstandalone_rtio_core_sed_selected328) | main_genericstandalone_rtio_core_sed_selected329) | main_genericstandalone_rtio_core_sed_selected330) | main_genericstandalone_rtio_core_sed_selected331) | main_genericstandalone_rtio_core_sed_selected332) | main_genericstandalone_rtio_core_sed_selected333) | main_genericstandalone_rtio_core_sed_selected334) | main_genericstandalone_rtio_core_sed_selected335);
	main_output_8x14_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected320 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected321 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected322 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected323 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected324 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected325 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected326 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected327 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected328 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected329 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected330 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected331 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected332 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected333 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected334 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected335 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x14_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected320 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected321 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected322 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected323 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected324 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected325 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected326 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected327 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected328 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected329 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected330 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected331 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected332 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected333 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected334 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected335 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x15_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected336 | main_genericstandalone_rtio_core_sed_selected337) | main_genericstandalone_rtio_core_sed_selected338) | main_genericstandalone_rtio_core_sed_selected339) | main_genericstandalone_rtio_core_sed_selected340) | main_genericstandalone_rtio_core_sed_selected341) | main_genericstandalone_rtio_core_sed_selected342) | main_genericstandalone_rtio_core_sed_selected343) | main_genericstandalone_rtio_core_sed_selected344) | main_genericstandalone_rtio_core_sed_selected345) | main_genericstandalone_rtio_core_sed_selected346) | main_genericstandalone_rtio_core_sed_selected347) | main_genericstandalone_rtio_core_sed_selected348) | main_genericstandalone_rtio_core_sed_selected349) | main_genericstandalone_rtio_core_sed_selected350) | main_genericstandalone_rtio_core_sed_selected351);
	main_output_8x15_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected336 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected337 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected338 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected339 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected340 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected341 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected342 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected343 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected344 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected345 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected346 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected347 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected348 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected349 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected350 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected351 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x15_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected336 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected337 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected338 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected339 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected340 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected341 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected342 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected343 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected344 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected345 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected346 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected347 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected348 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected349 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected350 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected351 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_spimaster1_ointerface1_stb0 <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected352 | main_genericstandalone_rtio_core_sed_selected353) | main_genericstandalone_rtio_core_sed_selected354) | main_genericstandalone_rtio_core_sed_selected355) | main_genericstandalone_rtio_core_sed_selected356) | main_genericstandalone_rtio_core_sed_selected357) | main_genericstandalone_rtio_core_sed_selected358) | main_genericstandalone_rtio_core_sed_selected359) | main_genericstandalone_rtio_core_sed_selected360) | main_genericstandalone_rtio_core_sed_selected361) | main_genericstandalone_rtio_core_sed_selected362) | main_genericstandalone_rtio_core_sed_selected363) | main_genericstandalone_rtio_core_sed_selected364) | main_genericstandalone_rtio_core_sed_selected365) | main_genericstandalone_rtio_core_sed_selected366) | main_genericstandalone_rtio_core_sed_selected367);
	main_spimaster1_ointerface1_address0 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected352 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected353 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected354 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected355 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected356 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected357 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected358 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected359 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected360 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected361 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected362 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected363 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected364 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected365 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected366 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected367 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_spimaster1_ointerface1_data0 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected352 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected353 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected354 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected355 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected356 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected357 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected358 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected359 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected360 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected361 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected362 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected363 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected364 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected365 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected366 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected367 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x1_stb1 <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected368 | main_genericstandalone_rtio_core_sed_selected369) | main_genericstandalone_rtio_core_sed_selected370) | main_genericstandalone_rtio_core_sed_selected371) | main_genericstandalone_rtio_core_sed_selected372) | main_genericstandalone_rtio_core_sed_selected373) | main_genericstandalone_rtio_core_sed_selected374) | main_genericstandalone_rtio_core_sed_selected375) | main_genericstandalone_rtio_core_sed_selected376) | main_genericstandalone_rtio_core_sed_selected377) | main_genericstandalone_rtio_core_sed_selected378) | main_genericstandalone_rtio_core_sed_selected379) | main_genericstandalone_rtio_core_sed_selected380) | main_genericstandalone_rtio_core_sed_selected381) | main_genericstandalone_rtio_core_sed_selected382) | main_genericstandalone_rtio_core_sed_selected383);
	main_output_8x1_fine_ts1 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected368 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected369 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected370 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected371 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected372 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected373 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected374 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected375 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected376 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected377 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected378 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected379 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected380 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected381 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected382 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected383 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x1_data1 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected368 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected369 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected370 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected371 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected372 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected373 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected374 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected375 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected376 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected377 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected378 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected379 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected380 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected381 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected382 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected383 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x16_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected384 | main_genericstandalone_rtio_core_sed_selected385) | main_genericstandalone_rtio_core_sed_selected386) | main_genericstandalone_rtio_core_sed_selected387) | main_genericstandalone_rtio_core_sed_selected388) | main_genericstandalone_rtio_core_sed_selected389) | main_genericstandalone_rtio_core_sed_selected390) | main_genericstandalone_rtio_core_sed_selected391) | main_genericstandalone_rtio_core_sed_selected392) | main_genericstandalone_rtio_core_sed_selected393) | main_genericstandalone_rtio_core_sed_selected394) | main_genericstandalone_rtio_core_sed_selected395) | main_genericstandalone_rtio_core_sed_selected396) | main_genericstandalone_rtio_core_sed_selected397) | main_genericstandalone_rtio_core_sed_selected398) | main_genericstandalone_rtio_core_sed_selected399);
	main_output_8x16_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected384 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected385 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected386 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected387 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected388 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected389 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected390 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected391 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected392 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected393 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected394 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected395 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected396 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected397 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected398 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected399 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x16_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected384 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected385 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected386 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected387 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected388 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected389 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected390 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected391 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected392 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected393 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected394 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected395 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected396 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected397 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected398 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected399 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x17_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected400 | main_genericstandalone_rtio_core_sed_selected401) | main_genericstandalone_rtio_core_sed_selected402) | main_genericstandalone_rtio_core_sed_selected403) | main_genericstandalone_rtio_core_sed_selected404) | main_genericstandalone_rtio_core_sed_selected405) | main_genericstandalone_rtio_core_sed_selected406) | main_genericstandalone_rtio_core_sed_selected407) | main_genericstandalone_rtio_core_sed_selected408) | main_genericstandalone_rtio_core_sed_selected409) | main_genericstandalone_rtio_core_sed_selected410) | main_genericstandalone_rtio_core_sed_selected411) | main_genericstandalone_rtio_core_sed_selected412) | main_genericstandalone_rtio_core_sed_selected413) | main_genericstandalone_rtio_core_sed_selected414) | main_genericstandalone_rtio_core_sed_selected415);
	main_output_8x17_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected400 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected401 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected402 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected403 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected404 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected405 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected406 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected407 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected408 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected409 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected410 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected411 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected412 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected413 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected414 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected415 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x17_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected400 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected401 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected402 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected403 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected404 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected405 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected406 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected407 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected408 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected409 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected410 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected411 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected412 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected413 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected414 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected415 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x18_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected416 | main_genericstandalone_rtio_core_sed_selected417) | main_genericstandalone_rtio_core_sed_selected418) | main_genericstandalone_rtio_core_sed_selected419) | main_genericstandalone_rtio_core_sed_selected420) | main_genericstandalone_rtio_core_sed_selected421) | main_genericstandalone_rtio_core_sed_selected422) | main_genericstandalone_rtio_core_sed_selected423) | main_genericstandalone_rtio_core_sed_selected424) | main_genericstandalone_rtio_core_sed_selected425) | main_genericstandalone_rtio_core_sed_selected426) | main_genericstandalone_rtio_core_sed_selected427) | main_genericstandalone_rtio_core_sed_selected428) | main_genericstandalone_rtio_core_sed_selected429) | main_genericstandalone_rtio_core_sed_selected430) | main_genericstandalone_rtio_core_sed_selected431);
	main_output_8x18_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected416 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected417 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected418 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected419 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected420 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected421 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected422 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected423 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected424 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected425 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected426 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected427 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected428 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected429 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected430 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected431 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x18_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected416 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected417 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected418 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected419 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected420 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected421 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected422 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected423 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected424 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected425 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected426 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected427 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected428 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected429 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected430 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected431 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x19_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected432 | main_genericstandalone_rtio_core_sed_selected433) | main_genericstandalone_rtio_core_sed_selected434) | main_genericstandalone_rtio_core_sed_selected435) | main_genericstandalone_rtio_core_sed_selected436) | main_genericstandalone_rtio_core_sed_selected437) | main_genericstandalone_rtio_core_sed_selected438) | main_genericstandalone_rtio_core_sed_selected439) | main_genericstandalone_rtio_core_sed_selected440) | main_genericstandalone_rtio_core_sed_selected441) | main_genericstandalone_rtio_core_sed_selected442) | main_genericstandalone_rtio_core_sed_selected443) | main_genericstandalone_rtio_core_sed_selected444) | main_genericstandalone_rtio_core_sed_selected445) | main_genericstandalone_rtio_core_sed_selected446) | main_genericstandalone_rtio_core_sed_selected447);
	main_output_8x19_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected432 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected433 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected434 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected435 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected436 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected437 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected438 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected439 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected440 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected441 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected442 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected443 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected444 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected445 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected446 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected447 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x19_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected432 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected433 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected434 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected435 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected436 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected437 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected438 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected439 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected440 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected441 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected442 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected443 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected444 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected445 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected446 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected447 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_spimaster0_ointerface0_stb1 <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected448 | main_genericstandalone_rtio_core_sed_selected449) | main_genericstandalone_rtio_core_sed_selected450) | main_genericstandalone_rtio_core_sed_selected451) | main_genericstandalone_rtio_core_sed_selected452) | main_genericstandalone_rtio_core_sed_selected453) | main_genericstandalone_rtio_core_sed_selected454) | main_genericstandalone_rtio_core_sed_selected455) | main_genericstandalone_rtio_core_sed_selected456) | main_genericstandalone_rtio_core_sed_selected457) | main_genericstandalone_rtio_core_sed_selected458) | main_genericstandalone_rtio_core_sed_selected459) | main_genericstandalone_rtio_core_sed_selected460) | main_genericstandalone_rtio_core_sed_selected461) | main_genericstandalone_rtio_core_sed_selected462) | main_genericstandalone_rtio_core_sed_selected463);
	main_spimaster0_ointerface0_address1 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected448 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected449 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected450 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected451 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected452 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected453 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected454 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected455 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected456 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected457 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected458 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected459 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected460 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected461 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected462 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected463 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_spimaster0_ointerface0_data1 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected448 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected449 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected450 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected451 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected452 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected453 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected454 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected455 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected456 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected457 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected458 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected459 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected460 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected461 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected462 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected463 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_spimaster1_ointerface1_stb1 <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected464 | main_genericstandalone_rtio_core_sed_selected465) | main_genericstandalone_rtio_core_sed_selected466) | main_genericstandalone_rtio_core_sed_selected467) | main_genericstandalone_rtio_core_sed_selected468) | main_genericstandalone_rtio_core_sed_selected469) | main_genericstandalone_rtio_core_sed_selected470) | main_genericstandalone_rtio_core_sed_selected471) | main_genericstandalone_rtio_core_sed_selected472) | main_genericstandalone_rtio_core_sed_selected473) | main_genericstandalone_rtio_core_sed_selected474) | main_genericstandalone_rtio_core_sed_selected475) | main_genericstandalone_rtio_core_sed_selected476) | main_genericstandalone_rtio_core_sed_selected477) | main_genericstandalone_rtio_core_sed_selected478) | main_genericstandalone_rtio_core_sed_selected479);
	main_spimaster1_ointerface1_address1 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected464 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected465 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected466 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected467 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected468 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected469 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected470 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected471 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected472 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected473 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected474 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected475 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected476 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected477 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected478 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected479 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_spimaster1_ointerface1_data1 <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected464 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected465 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected466 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected467 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected468 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected469 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected470 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected471 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected472 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected473 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected474 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected475 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected476 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected477 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected478 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected479 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output_8x20_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected480 | main_genericstandalone_rtio_core_sed_selected481) | main_genericstandalone_rtio_core_sed_selected482) | main_genericstandalone_rtio_core_sed_selected483) | main_genericstandalone_rtio_core_sed_selected484) | main_genericstandalone_rtio_core_sed_selected485) | main_genericstandalone_rtio_core_sed_selected486) | main_genericstandalone_rtio_core_sed_selected487) | main_genericstandalone_rtio_core_sed_selected488) | main_genericstandalone_rtio_core_sed_selected489) | main_genericstandalone_rtio_core_sed_selected490) | main_genericstandalone_rtio_core_sed_selected491) | main_genericstandalone_rtio_core_sed_selected492) | main_genericstandalone_rtio_core_sed_selected493) | main_genericstandalone_rtio_core_sed_selected494) | main_genericstandalone_rtio_core_sed_selected495);
	main_output_8x20_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected480 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected481 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected482 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected483 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected484 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected485 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected486 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected487 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected488 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected489 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected490 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected491 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected492 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected493 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected494 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected495 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x20_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected480 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected481 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected482 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected483 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected484 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected485 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected486 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected487 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected488 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected489 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected490 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected491 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected492 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected493 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected494 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected495 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_spimaster2_ointerface2_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected496 | main_genericstandalone_rtio_core_sed_selected497) | main_genericstandalone_rtio_core_sed_selected498) | main_genericstandalone_rtio_core_sed_selected499) | main_genericstandalone_rtio_core_sed_selected500) | main_genericstandalone_rtio_core_sed_selected501) | main_genericstandalone_rtio_core_sed_selected502) | main_genericstandalone_rtio_core_sed_selected503) | main_genericstandalone_rtio_core_sed_selected504) | main_genericstandalone_rtio_core_sed_selected505) | main_genericstandalone_rtio_core_sed_selected506) | main_genericstandalone_rtio_core_sed_selected507) | main_genericstandalone_rtio_core_sed_selected508) | main_genericstandalone_rtio_core_sed_selected509) | main_genericstandalone_rtio_core_sed_selected510) | main_genericstandalone_rtio_core_sed_selected511);
	main_spimaster2_ointerface2_address <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected496 ? main_genericstandalone_rtio_core_sed_record0_payload_address2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected497 ? main_genericstandalone_rtio_core_sed_record1_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected498 ? main_genericstandalone_rtio_core_sed_record2_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected499 ? main_genericstandalone_rtio_core_sed_record3_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected500 ? main_genericstandalone_rtio_core_sed_record4_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected501 ? main_genericstandalone_rtio_core_sed_record5_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected502 ? main_genericstandalone_rtio_core_sed_record6_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected503 ? main_genericstandalone_rtio_core_sed_record7_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected504 ? main_genericstandalone_rtio_core_sed_record8_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected505 ? main_genericstandalone_rtio_core_sed_record9_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected506 ? main_genericstandalone_rtio_core_sed_record10_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected507 ? main_genericstandalone_rtio_core_sed_record11_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected508 ? main_genericstandalone_rtio_core_sed_record12_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected509 ? main_genericstandalone_rtio_core_sed_record13_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected510 ? main_genericstandalone_rtio_core_sed_record14_payload_address2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected511 ? main_genericstandalone_rtio_core_sed_record15_payload_address2 : 1'd0));
	main_spimaster2_ointerface2_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected496 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected497 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected498 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected499 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected500 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected501 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected502 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected503 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected504 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected505 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected506 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected507 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected508 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected509 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected510 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected511 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_ldac_phy_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected512 | main_genericstandalone_rtio_core_sed_selected513) | main_genericstandalone_rtio_core_sed_selected514) | main_genericstandalone_rtio_core_sed_selected515) | main_genericstandalone_rtio_core_sed_selected516) | main_genericstandalone_rtio_core_sed_selected517) | main_genericstandalone_rtio_core_sed_selected518) | main_genericstandalone_rtio_core_sed_selected519) | main_genericstandalone_rtio_core_sed_selected520) | main_genericstandalone_rtio_core_sed_selected521) | main_genericstandalone_rtio_core_sed_selected522) | main_genericstandalone_rtio_core_sed_selected523) | main_genericstandalone_rtio_core_sed_selected524) | main_genericstandalone_rtio_core_sed_selected525) | main_genericstandalone_rtio_core_sed_selected526) | main_genericstandalone_rtio_core_sed_selected527);
	main_ldac_phy_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected512 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected513 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected514 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected515 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected516 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected517 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected518 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected519 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected520 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected521 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected522 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected523 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected524 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected525 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected526 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected527 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_ldac_phy_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected512 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected513 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected514 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected515 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected516 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected517 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected518 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected519 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected520 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected521 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected522 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected523 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected524 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected525 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected526 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected527 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_clr_phy_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected528 | main_genericstandalone_rtio_core_sed_selected529) | main_genericstandalone_rtio_core_sed_selected530) | main_genericstandalone_rtio_core_sed_selected531) | main_genericstandalone_rtio_core_sed_selected532) | main_genericstandalone_rtio_core_sed_selected533) | main_genericstandalone_rtio_core_sed_selected534) | main_genericstandalone_rtio_core_sed_selected535) | main_genericstandalone_rtio_core_sed_selected536) | main_genericstandalone_rtio_core_sed_selected537) | main_genericstandalone_rtio_core_sed_selected538) | main_genericstandalone_rtio_core_sed_selected539) | main_genericstandalone_rtio_core_sed_selected540) | main_genericstandalone_rtio_core_sed_selected541) | main_genericstandalone_rtio_core_sed_selected542) | main_genericstandalone_rtio_core_sed_selected543);
	main_clr_phy_fine_ts <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected528 ? main_genericstandalone_rtio_core_sed_record0_payload_fine_ts1[2:0] : 1'd0) | (main_genericstandalone_rtio_core_sed_selected529 ? main_genericstandalone_rtio_core_sed_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected530 ? main_genericstandalone_rtio_core_sed_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected531 ? main_genericstandalone_rtio_core_sed_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected532 ? main_genericstandalone_rtio_core_sed_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected533 ? main_genericstandalone_rtio_core_sed_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected534 ? main_genericstandalone_rtio_core_sed_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected535 ? main_genericstandalone_rtio_core_sed_record7_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected536 ? main_genericstandalone_rtio_core_sed_record8_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected537 ? main_genericstandalone_rtio_core_sed_record9_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected538 ? main_genericstandalone_rtio_core_sed_record10_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected539 ? main_genericstandalone_rtio_core_sed_record11_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected540 ? main_genericstandalone_rtio_core_sed_record12_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected541 ? main_genericstandalone_rtio_core_sed_record13_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected542 ? main_genericstandalone_rtio_core_sed_record14_payload_fine_ts1[2:0] : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected543 ? main_genericstandalone_rtio_core_sed_record15_payload_fine_ts1[2:0] : 1'd0));
	main_clr_phy_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected528 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected529 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected530 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected531 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected532 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected533 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected534 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected535 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected536 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected537 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected538 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected539 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected540 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected541 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected542 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected543 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output0_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected544 | main_genericstandalone_rtio_core_sed_selected545) | main_genericstandalone_rtio_core_sed_selected546) | main_genericstandalone_rtio_core_sed_selected547) | main_genericstandalone_rtio_core_sed_selected548) | main_genericstandalone_rtio_core_sed_selected549) | main_genericstandalone_rtio_core_sed_selected550) | main_genericstandalone_rtio_core_sed_selected551) | main_genericstandalone_rtio_core_sed_selected552) | main_genericstandalone_rtio_core_sed_selected553) | main_genericstandalone_rtio_core_sed_selected554) | main_genericstandalone_rtio_core_sed_selected555) | main_genericstandalone_rtio_core_sed_selected556) | main_genericstandalone_rtio_core_sed_selected557) | main_genericstandalone_rtio_core_sed_selected558) | main_genericstandalone_rtio_core_sed_selected559);
	main_output0_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected544 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected545 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected546 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected547 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected548 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected549 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected550 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected551 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected552 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected553 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected554 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected555 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected556 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected557 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected558 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected559 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output1_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected560 | main_genericstandalone_rtio_core_sed_selected561) | main_genericstandalone_rtio_core_sed_selected562) | main_genericstandalone_rtio_core_sed_selected563) | main_genericstandalone_rtio_core_sed_selected564) | main_genericstandalone_rtio_core_sed_selected565) | main_genericstandalone_rtio_core_sed_selected566) | main_genericstandalone_rtio_core_sed_selected567) | main_genericstandalone_rtio_core_sed_selected568) | main_genericstandalone_rtio_core_sed_selected569) | main_genericstandalone_rtio_core_sed_selected570) | main_genericstandalone_rtio_core_sed_selected571) | main_genericstandalone_rtio_core_sed_selected572) | main_genericstandalone_rtio_core_sed_selected573) | main_genericstandalone_rtio_core_sed_selected574) | main_genericstandalone_rtio_core_sed_selected575);
	main_output1_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected560 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected561 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected562 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected563 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected564 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected565 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected566 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected567 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected568 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected569 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected570 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected571 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected572 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected573 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected574 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected575 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_output2_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected576 | main_genericstandalone_rtio_core_sed_selected577) | main_genericstandalone_rtio_core_sed_selected578) | main_genericstandalone_rtio_core_sed_selected579) | main_genericstandalone_rtio_core_sed_selected580) | main_genericstandalone_rtio_core_sed_selected581) | main_genericstandalone_rtio_core_sed_selected582) | main_genericstandalone_rtio_core_sed_selected583) | main_genericstandalone_rtio_core_sed_selected584) | main_genericstandalone_rtio_core_sed_selected585) | main_genericstandalone_rtio_core_sed_selected586) | main_genericstandalone_rtio_core_sed_selected587) | main_genericstandalone_rtio_core_sed_selected588) | main_genericstandalone_rtio_core_sed_selected589) | main_genericstandalone_rtio_core_sed_selected590) | main_genericstandalone_rtio_core_sed_selected591);
	main_output2_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected576 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected577 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected578 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected579 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected580 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected581 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected582 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected583 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected584 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected585 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected586 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected587 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected588 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected589 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected590 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected591 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_stb <= (((((((((((((((main_genericstandalone_rtio_core_sed_selected592 | main_genericstandalone_rtio_core_sed_selected593) | main_genericstandalone_rtio_core_sed_selected594) | main_genericstandalone_rtio_core_sed_selected595) | main_genericstandalone_rtio_core_sed_selected596) | main_genericstandalone_rtio_core_sed_selected597) | main_genericstandalone_rtio_core_sed_selected598) | main_genericstandalone_rtio_core_sed_selected599) | main_genericstandalone_rtio_core_sed_selected600) | main_genericstandalone_rtio_core_sed_selected601) | main_genericstandalone_rtio_core_sed_selected602) | main_genericstandalone_rtio_core_sed_selected603) | main_genericstandalone_rtio_core_sed_selected604) | main_genericstandalone_rtio_core_sed_selected605) | main_genericstandalone_rtio_core_sed_selected606) | main_genericstandalone_rtio_core_sed_selected607);
	main_data <= ((((((((((((((((main_genericstandalone_rtio_core_sed_selected592 ? main_genericstandalone_rtio_core_sed_record0_payload_data2 : 1'd0) | (main_genericstandalone_rtio_core_sed_selected593 ? main_genericstandalone_rtio_core_sed_record1_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected594 ? main_genericstandalone_rtio_core_sed_record2_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected595 ? main_genericstandalone_rtio_core_sed_record3_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected596 ? main_genericstandalone_rtio_core_sed_record4_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected597 ? main_genericstandalone_rtio_core_sed_record5_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected598 ? main_genericstandalone_rtio_core_sed_record6_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected599 ? main_genericstandalone_rtio_core_sed_record7_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected600 ? main_genericstandalone_rtio_core_sed_record8_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected601 ? main_genericstandalone_rtio_core_sed_record9_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected602 ? main_genericstandalone_rtio_core_sed_record10_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected603 ? main_genericstandalone_rtio_core_sed_record11_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected604 ? main_genericstandalone_rtio_core_sed_record12_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected605 ? main_genericstandalone_rtio_core_sed_record13_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected606 ? main_genericstandalone_rtio_core_sed_record14_payload_data2 : 1'd0)) | (main_genericstandalone_rtio_core_sed_selected607 ? main_genericstandalone_rtio_core_sed_record15_payload_data2 : 1'd0));
	main_genericstandalone_rtio_core_sed_busy <= 1'd0;
	main_genericstandalone_rtio_core_sed_busy_channel <= 1'd0;
	main_genericstandalone_rtio_core_sed_stb_r0 <= (main_genericstandalone_rtio_core_sed_record0_valid1 & (~main_genericstandalone_rtio_core_sed_record0_collision));
	main_genericstandalone_rtio_core_sed_channel_r0 <= main_genericstandalone_rtio_core_sed_record0_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r0 & builder_sync_basiclowerer_self0)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r0;
	end
	main_genericstandalone_rtio_core_sed_stb_r1 <= (main_genericstandalone_rtio_core_sed_record1_valid1 & (~main_genericstandalone_rtio_core_sed_record1_collision));
	main_genericstandalone_rtio_core_sed_channel_r1 <= main_genericstandalone_rtio_core_sed_record1_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r1 & builder_sync_basiclowerer_self1)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r1;
	end
	main_genericstandalone_rtio_core_sed_stb_r2 <= (main_genericstandalone_rtio_core_sed_record2_valid1 & (~main_genericstandalone_rtio_core_sed_record2_collision));
	main_genericstandalone_rtio_core_sed_channel_r2 <= main_genericstandalone_rtio_core_sed_record2_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r2 & builder_sync_basiclowerer_self2)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r2;
	end
	main_genericstandalone_rtio_core_sed_stb_r3 <= (main_genericstandalone_rtio_core_sed_record3_valid1 & (~main_genericstandalone_rtio_core_sed_record3_collision));
	main_genericstandalone_rtio_core_sed_channel_r3 <= main_genericstandalone_rtio_core_sed_record3_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r3 & builder_sync_basiclowerer_self3)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r3;
	end
	main_genericstandalone_rtio_core_sed_stb_r4 <= (main_genericstandalone_rtio_core_sed_record4_valid1 & (~main_genericstandalone_rtio_core_sed_record4_collision));
	main_genericstandalone_rtio_core_sed_channel_r4 <= main_genericstandalone_rtio_core_sed_record4_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r4 & builder_sync_basiclowerer_self4)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r4;
	end
	main_genericstandalone_rtio_core_sed_stb_r5 <= (main_genericstandalone_rtio_core_sed_record5_valid1 & (~main_genericstandalone_rtio_core_sed_record5_collision));
	main_genericstandalone_rtio_core_sed_channel_r5 <= main_genericstandalone_rtio_core_sed_record5_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r5 & builder_sync_basiclowerer_self5)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r5;
	end
	main_genericstandalone_rtio_core_sed_stb_r6 <= (main_genericstandalone_rtio_core_sed_record6_valid1 & (~main_genericstandalone_rtio_core_sed_record6_collision));
	main_genericstandalone_rtio_core_sed_channel_r6 <= main_genericstandalone_rtio_core_sed_record6_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r6 & builder_sync_basiclowerer_self6)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r6;
	end
	main_genericstandalone_rtio_core_sed_stb_r7 <= (main_genericstandalone_rtio_core_sed_record7_valid1 & (~main_genericstandalone_rtio_core_sed_record7_collision));
	main_genericstandalone_rtio_core_sed_channel_r7 <= main_genericstandalone_rtio_core_sed_record7_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r7 & builder_sync_basiclowerer_self7)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r7;
	end
	main_genericstandalone_rtio_core_sed_stb_r8 <= (main_genericstandalone_rtio_core_sed_record8_valid1 & (~main_genericstandalone_rtio_core_sed_record8_collision));
	main_genericstandalone_rtio_core_sed_channel_r8 <= main_genericstandalone_rtio_core_sed_record8_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r8 & builder_sync_basiclowerer_self8)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r8;
	end
	main_genericstandalone_rtio_core_sed_stb_r9 <= (main_genericstandalone_rtio_core_sed_record9_valid1 & (~main_genericstandalone_rtio_core_sed_record9_collision));
	main_genericstandalone_rtio_core_sed_channel_r9 <= main_genericstandalone_rtio_core_sed_record9_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r9 & builder_sync_basiclowerer_self9)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r9;
	end
	main_genericstandalone_rtio_core_sed_stb_r10 <= (main_genericstandalone_rtio_core_sed_record10_valid1 & (~main_genericstandalone_rtio_core_sed_record10_collision));
	main_genericstandalone_rtio_core_sed_channel_r10 <= main_genericstandalone_rtio_core_sed_record10_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r10 & builder_sync_basiclowerer_self10)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r10;
	end
	main_genericstandalone_rtio_core_sed_stb_r11 <= (main_genericstandalone_rtio_core_sed_record11_valid1 & (~main_genericstandalone_rtio_core_sed_record11_collision));
	main_genericstandalone_rtio_core_sed_channel_r11 <= main_genericstandalone_rtio_core_sed_record11_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r11 & builder_sync_basiclowerer_self11)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r11;
	end
	main_genericstandalone_rtio_core_sed_stb_r12 <= (main_genericstandalone_rtio_core_sed_record12_valid1 & (~main_genericstandalone_rtio_core_sed_record12_collision));
	main_genericstandalone_rtio_core_sed_channel_r12 <= main_genericstandalone_rtio_core_sed_record12_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r12 & builder_sync_basiclowerer_self12)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r12;
	end
	main_genericstandalone_rtio_core_sed_stb_r13 <= (main_genericstandalone_rtio_core_sed_record13_valid1 & (~main_genericstandalone_rtio_core_sed_record13_collision));
	main_genericstandalone_rtio_core_sed_channel_r13 <= main_genericstandalone_rtio_core_sed_record13_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r13 & builder_sync_basiclowerer_self13)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r13;
	end
	main_genericstandalone_rtio_core_sed_stb_r14 <= (main_genericstandalone_rtio_core_sed_record14_valid1 & (~main_genericstandalone_rtio_core_sed_record14_collision));
	main_genericstandalone_rtio_core_sed_channel_r14 <= main_genericstandalone_rtio_core_sed_record14_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r14 & builder_sync_basiclowerer_self14)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r14;
	end
	main_genericstandalone_rtio_core_sed_stb_r15 <= (main_genericstandalone_rtio_core_sed_record15_valid1 & (~main_genericstandalone_rtio_core_sed_record15_collision));
	main_genericstandalone_rtio_core_sed_channel_r15 <= main_genericstandalone_rtio_core_sed_record15_payload_channel2;
	if ((main_genericstandalone_rtio_core_sed_stb_r15 & builder_sync_basiclowerer_self15)) begin
		main_genericstandalone_rtio_core_sed_busy <= 1'd1;
		main_genericstandalone_rtio_core_sed_busy_channel <= main_genericstandalone_rtio_core_sed_channel_r15;
	end
	if (({(~main_genericstandalone_rtio_core_sed_record0_valid0), main_genericstandalone_rtio_core_sed_record0_payload_channel1} == {(~main_genericstandalone_rtio_core_sed_record1_valid0), main_genericstandalone_rtio_core_sed_record1_payload_channel1})) begin
		if (((((main_genericstandalone_rtio_core_sed_record0_seqn1[11] == main_genericstandalone_rtio_core_sed_record0_seqn1[12]) & (main_genericstandalone_rtio_core_sed_record1_seqn1[11] == main_genericstandalone_rtio_core_sed_record1_seqn1[12])) & (main_genericstandalone_rtio_core_sed_record0_seqn1[12] != main_genericstandalone_rtio_core_sed_record1_seqn1[12])) ? main_genericstandalone_rtio_core_sed_record0_seqn1[12] : (main_genericstandalone_rtio_core_sed_record0_seqn1 < main_genericstandalone_rtio_core_sed_record1_seqn1))) begin
			main_genericstandalone_rtio_core_sed_record0_rec_valid <= main_genericstandalone_rtio_core_sed_record1_valid0;
			main_genericstandalone_rtio_core_sed_record0_rec_seqn <= main_genericstandalone_rtio_core_sed_record1_seqn1;
			main_genericstandalone_rtio_core_sed_record0_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record1_replace_occured;
			main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record1_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record1_payload_channel1;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record1_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_address <= main_genericstandalone_rtio_core_sed_record1_payload_address1;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_data <= main_genericstandalone_rtio_core_sed_record1_payload_data1;
			main_genericstandalone_rtio_core_sed_record1_rec_valid <= main_genericstandalone_rtio_core_sed_record0_valid0;
			main_genericstandalone_rtio_core_sed_record1_rec_seqn <= main_genericstandalone_rtio_core_sed_record0_seqn1;
			main_genericstandalone_rtio_core_sed_record1_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record0_replace_occured;
			main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record0_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record0_payload_channel1;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record0_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_address <= main_genericstandalone_rtio_core_sed_record0_payload_address1;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_data <= main_genericstandalone_rtio_core_sed_record0_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record0_rec_valid <= main_genericstandalone_rtio_core_sed_record0_valid0;
			main_genericstandalone_rtio_core_sed_record0_rec_seqn <= main_genericstandalone_rtio_core_sed_record0_seqn1;
			main_genericstandalone_rtio_core_sed_record0_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record0_replace_occured;
			main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record0_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record0_payload_channel1;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record0_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_address <= main_genericstandalone_rtio_core_sed_record0_payload_address1;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_data <= main_genericstandalone_rtio_core_sed_record0_payload_data1;
			main_genericstandalone_rtio_core_sed_record1_rec_valid <= main_genericstandalone_rtio_core_sed_record1_valid0;
			main_genericstandalone_rtio_core_sed_record1_rec_seqn <= main_genericstandalone_rtio_core_sed_record1_seqn1;
			main_genericstandalone_rtio_core_sed_record1_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record1_replace_occured;
			main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record1_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record1_payload_channel1;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record1_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_address <= main_genericstandalone_rtio_core_sed_record1_payload_address1;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_data <= main_genericstandalone_rtio_core_sed_record1_payload_data1;
		end
		main_genericstandalone_rtio_core_sed_record0_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference0;
		main_genericstandalone_rtio_core_sed_record1_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record0_valid0), main_genericstandalone_rtio_core_sed_record0_payload_channel1} < {(~main_genericstandalone_rtio_core_sed_record1_valid0), main_genericstandalone_rtio_core_sed_record1_payload_channel1})) begin
			main_genericstandalone_rtio_core_sed_record0_rec_valid <= main_genericstandalone_rtio_core_sed_record0_valid0;
			main_genericstandalone_rtio_core_sed_record0_rec_seqn <= main_genericstandalone_rtio_core_sed_record0_seqn1;
			main_genericstandalone_rtio_core_sed_record0_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record0_replace_occured;
			main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record0_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record0_payload_channel1;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record0_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_address <= main_genericstandalone_rtio_core_sed_record0_payload_address1;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_data <= main_genericstandalone_rtio_core_sed_record0_payload_data1;
			main_genericstandalone_rtio_core_sed_record1_rec_valid <= main_genericstandalone_rtio_core_sed_record1_valid0;
			main_genericstandalone_rtio_core_sed_record1_rec_seqn <= main_genericstandalone_rtio_core_sed_record1_seqn1;
			main_genericstandalone_rtio_core_sed_record1_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record1_replace_occured;
			main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record1_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record1_payload_channel1;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record1_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_address <= main_genericstandalone_rtio_core_sed_record1_payload_address1;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_data <= main_genericstandalone_rtio_core_sed_record1_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record0_rec_valid <= main_genericstandalone_rtio_core_sed_record1_valid0;
			main_genericstandalone_rtio_core_sed_record0_rec_seqn <= main_genericstandalone_rtio_core_sed_record1_seqn1;
			main_genericstandalone_rtio_core_sed_record0_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record1_replace_occured;
			main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record1_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record1_payload_channel1;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record1_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_address <= main_genericstandalone_rtio_core_sed_record1_payload_address1;
			main_genericstandalone_rtio_core_sed_record0_rec_payload_data <= main_genericstandalone_rtio_core_sed_record1_payload_data1;
			main_genericstandalone_rtio_core_sed_record1_rec_valid <= main_genericstandalone_rtio_core_sed_record0_valid0;
			main_genericstandalone_rtio_core_sed_record1_rec_seqn <= main_genericstandalone_rtio_core_sed_record0_seqn1;
			main_genericstandalone_rtio_core_sed_record1_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record0_replace_occured;
			main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record0_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record0_payload_channel1;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record0_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_address <= main_genericstandalone_rtio_core_sed_record0_payload_address1;
			main_genericstandalone_rtio_core_sed_record1_rec_payload_data <= main_genericstandalone_rtio_core_sed_record0_payload_data1;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record2_valid0), main_genericstandalone_rtio_core_sed_record2_payload_channel1} == {(~main_genericstandalone_rtio_core_sed_record3_valid0), main_genericstandalone_rtio_core_sed_record3_payload_channel1})) begin
		if (((((main_genericstandalone_rtio_core_sed_record2_seqn1[11] == main_genericstandalone_rtio_core_sed_record2_seqn1[12]) & (main_genericstandalone_rtio_core_sed_record3_seqn1[11] == main_genericstandalone_rtio_core_sed_record3_seqn1[12])) & (main_genericstandalone_rtio_core_sed_record2_seqn1[12] != main_genericstandalone_rtio_core_sed_record3_seqn1[12])) ? main_genericstandalone_rtio_core_sed_record2_seqn1[12] : (main_genericstandalone_rtio_core_sed_record2_seqn1 < main_genericstandalone_rtio_core_sed_record3_seqn1))) begin
			main_genericstandalone_rtio_core_sed_record2_rec_valid <= main_genericstandalone_rtio_core_sed_record3_valid0;
			main_genericstandalone_rtio_core_sed_record2_rec_seqn <= main_genericstandalone_rtio_core_sed_record3_seqn1;
			main_genericstandalone_rtio_core_sed_record2_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record3_replace_occured;
			main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record3_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record3_payload_channel1;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record3_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_address <= main_genericstandalone_rtio_core_sed_record3_payload_address1;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_data <= main_genericstandalone_rtio_core_sed_record3_payload_data1;
			main_genericstandalone_rtio_core_sed_record3_rec_valid <= main_genericstandalone_rtio_core_sed_record2_valid0;
			main_genericstandalone_rtio_core_sed_record3_rec_seqn <= main_genericstandalone_rtio_core_sed_record2_seqn1;
			main_genericstandalone_rtio_core_sed_record3_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record2_replace_occured;
			main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record2_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record2_payload_channel1;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record2_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_address <= main_genericstandalone_rtio_core_sed_record2_payload_address1;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_data <= main_genericstandalone_rtio_core_sed_record2_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record2_rec_valid <= main_genericstandalone_rtio_core_sed_record2_valid0;
			main_genericstandalone_rtio_core_sed_record2_rec_seqn <= main_genericstandalone_rtio_core_sed_record2_seqn1;
			main_genericstandalone_rtio_core_sed_record2_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record2_replace_occured;
			main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record2_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record2_payload_channel1;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record2_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_address <= main_genericstandalone_rtio_core_sed_record2_payload_address1;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_data <= main_genericstandalone_rtio_core_sed_record2_payload_data1;
			main_genericstandalone_rtio_core_sed_record3_rec_valid <= main_genericstandalone_rtio_core_sed_record3_valid0;
			main_genericstandalone_rtio_core_sed_record3_rec_seqn <= main_genericstandalone_rtio_core_sed_record3_seqn1;
			main_genericstandalone_rtio_core_sed_record3_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record3_replace_occured;
			main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record3_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record3_payload_channel1;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record3_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_address <= main_genericstandalone_rtio_core_sed_record3_payload_address1;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_data <= main_genericstandalone_rtio_core_sed_record3_payload_data1;
		end
		main_genericstandalone_rtio_core_sed_record2_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference1;
		main_genericstandalone_rtio_core_sed_record3_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record2_valid0), main_genericstandalone_rtio_core_sed_record2_payload_channel1} < {(~main_genericstandalone_rtio_core_sed_record3_valid0), main_genericstandalone_rtio_core_sed_record3_payload_channel1})) begin
			main_genericstandalone_rtio_core_sed_record2_rec_valid <= main_genericstandalone_rtio_core_sed_record2_valid0;
			main_genericstandalone_rtio_core_sed_record2_rec_seqn <= main_genericstandalone_rtio_core_sed_record2_seqn1;
			main_genericstandalone_rtio_core_sed_record2_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record2_replace_occured;
			main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record2_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record2_payload_channel1;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record2_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_address <= main_genericstandalone_rtio_core_sed_record2_payload_address1;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_data <= main_genericstandalone_rtio_core_sed_record2_payload_data1;
			main_genericstandalone_rtio_core_sed_record3_rec_valid <= main_genericstandalone_rtio_core_sed_record3_valid0;
			main_genericstandalone_rtio_core_sed_record3_rec_seqn <= main_genericstandalone_rtio_core_sed_record3_seqn1;
			main_genericstandalone_rtio_core_sed_record3_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record3_replace_occured;
			main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record3_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record3_payload_channel1;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record3_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_address <= main_genericstandalone_rtio_core_sed_record3_payload_address1;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_data <= main_genericstandalone_rtio_core_sed_record3_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record2_rec_valid <= main_genericstandalone_rtio_core_sed_record3_valid0;
			main_genericstandalone_rtio_core_sed_record2_rec_seqn <= main_genericstandalone_rtio_core_sed_record3_seqn1;
			main_genericstandalone_rtio_core_sed_record2_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record3_replace_occured;
			main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record3_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record3_payload_channel1;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record3_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_address <= main_genericstandalone_rtio_core_sed_record3_payload_address1;
			main_genericstandalone_rtio_core_sed_record2_rec_payload_data <= main_genericstandalone_rtio_core_sed_record3_payload_data1;
			main_genericstandalone_rtio_core_sed_record3_rec_valid <= main_genericstandalone_rtio_core_sed_record2_valid0;
			main_genericstandalone_rtio_core_sed_record3_rec_seqn <= main_genericstandalone_rtio_core_sed_record2_seqn1;
			main_genericstandalone_rtio_core_sed_record3_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record2_replace_occured;
			main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record2_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record2_payload_channel1;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record2_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_address <= main_genericstandalone_rtio_core_sed_record2_payload_address1;
			main_genericstandalone_rtio_core_sed_record3_rec_payload_data <= main_genericstandalone_rtio_core_sed_record2_payload_data1;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record4_valid0), main_genericstandalone_rtio_core_sed_record4_payload_channel1} == {(~main_genericstandalone_rtio_core_sed_record5_valid0), main_genericstandalone_rtio_core_sed_record5_payload_channel1})) begin
		if (((((main_genericstandalone_rtio_core_sed_record4_seqn1[11] == main_genericstandalone_rtio_core_sed_record4_seqn1[12]) & (main_genericstandalone_rtio_core_sed_record5_seqn1[11] == main_genericstandalone_rtio_core_sed_record5_seqn1[12])) & (main_genericstandalone_rtio_core_sed_record4_seqn1[12] != main_genericstandalone_rtio_core_sed_record5_seqn1[12])) ? main_genericstandalone_rtio_core_sed_record4_seqn1[12] : (main_genericstandalone_rtio_core_sed_record4_seqn1 < main_genericstandalone_rtio_core_sed_record5_seqn1))) begin
			main_genericstandalone_rtio_core_sed_record4_rec_valid <= main_genericstandalone_rtio_core_sed_record5_valid0;
			main_genericstandalone_rtio_core_sed_record4_rec_seqn <= main_genericstandalone_rtio_core_sed_record5_seqn1;
			main_genericstandalone_rtio_core_sed_record4_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record5_replace_occured;
			main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record5_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record5_payload_channel1;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record5_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_address <= main_genericstandalone_rtio_core_sed_record5_payload_address1;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_data <= main_genericstandalone_rtio_core_sed_record5_payload_data1;
			main_genericstandalone_rtio_core_sed_record5_rec_valid <= main_genericstandalone_rtio_core_sed_record4_valid0;
			main_genericstandalone_rtio_core_sed_record5_rec_seqn <= main_genericstandalone_rtio_core_sed_record4_seqn1;
			main_genericstandalone_rtio_core_sed_record5_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record4_replace_occured;
			main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record4_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record4_payload_channel1;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record4_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_address <= main_genericstandalone_rtio_core_sed_record4_payload_address1;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_data <= main_genericstandalone_rtio_core_sed_record4_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record4_rec_valid <= main_genericstandalone_rtio_core_sed_record4_valid0;
			main_genericstandalone_rtio_core_sed_record4_rec_seqn <= main_genericstandalone_rtio_core_sed_record4_seqn1;
			main_genericstandalone_rtio_core_sed_record4_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record4_replace_occured;
			main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record4_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record4_payload_channel1;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record4_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_address <= main_genericstandalone_rtio_core_sed_record4_payload_address1;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_data <= main_genericstandalone_rtio_core_sed_record4_payload_data1;
			main_genericstandalone_rtio_core_sed_record5_rec_valid <= main_genericstandalone_rtio_core_sed_record5_valid0;
			main_genericstandalone_rtio_core_sed_record5_rec_seqn <= main_genericstandalone_rtio_core_sed_record5_seqn1;
			main_genericstandalone_rtio_core_sed_record5_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record5_replace_occured;
			main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record5_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record5_payload_channel1;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record5_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_address <= main_genericstandalone_rtio_core_sed_record5_payload_address1;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_data <= main_genericstandalone_rtio_core_sed_record5_payload_data1;
		end
		main_genericstandalone_rtio_core_sed_record4_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference2;
		main_genericstandalone_rtio_core_sed_record5_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record4_valid0), main_genericstandalone_rtio_core_sed_record4_payload_channel1} < {(~main_genericstandalone_rtio_core_sed_record5_valid0), main_genericstandalone_rtio_core_sed_record5_payload_channel1})) begin
			main_genericstandalone_rtio_core_sed_record4_rec_valid <= main_genericstandalone_rtio_core_sed_record4_valid0;
			main_genericstandalone_rtio_core_sed_record4_rec_seqn <= main_genericstandalone_rtio_core_sed_record4_seqn1;
			main_genericstandalone_rtio_core_sed_record4_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record4_replace_occured;
			main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record4_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record4_payload_channel1;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record4_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_address <= main_genericstandalone_rtio_core_sed_record4_payload_address1;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_data <= main_genericstandalone_rtio_core_sed_record4_payload_data1;
			main_genericstandalone_rtio_core_sed_record5_rec_valid <= main_genericstandalone_rtio_core_sed_record5_valid0;
			main_genericstandalone_rtio_core_sed_record5_rec_seqn <= main_genericstandalone_rtio_core_sed_record5_seqn1;
			main_genericstandalone_rtio_core_sed_record5_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record5_replace_occured;
			main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record5_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record5_payload_channel1;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record5_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_address <= main_genericstandalone_rtio_core_sed_record5_payload_address1;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_data <= main_genericstandalone_rtio_core_sed_record5_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record4_rec_valid <= main_genericstandalone_rtio_core_sed_record5_valid0;
			main_genericstandalone_rtio_core_sed_record4_rec_seqn <= main_genericstandalone_rtio_core_sed_record5_seqn1;
			main_genericstandalone_rtio_core_sed_record4_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record5_replace_occured;
			main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record5_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record5_payload_channel1;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record5_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_address <= main_genericstandalone_rtio_core_sed_record5_payload_address1;
			main_genericstandalone_rtio_core_sed_record4_rec_payload_data <= main_genericstandalone_rtio_core_sed_record5_payload_data1;
			main_genericstandalone_rtio_core_sed_record5_rec_valid <= main_genericstandalone_rtio_core_sed_record4_valid0;
			main_genericstandalone_rtio_core_sed_record5_rec_seqn <= main_genericstandalone_rtio_core_sed_record4_seqn1;
			main_genericstandalone_rtio_core_sed_record5_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record4_replace_occured;
			main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record4_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record4_payload_channel1;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record4_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_address <= main_genericstandalone_rtio_core_sed_record4_payload_address1;
			main_genericstandalone_rtio_core_sed_record5_rec_payload_data <= main_genericstandalone_rtio_core_sed_record4_payload_data1;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record6_valid0), main_genericstandalone_rtio_core_sed_record6_payload_channel1} == {(~main_genericstandalone_rtio_core_sed_record7_valid0), main_genericstandalone_rtio_core_sed_record7_payload_channel1})) begin
		if (((((main_genericstandalone_rtio_core_sed_record6_seqn1[11] == main_genericstandalone_rtio_core_sed_record6_seqn1[12]) & (main_genericstandalone_rtio_core_sed_record7_seqn1[11] == main_genericstandalone_rtio_core_sed_record7_seqn1[12])) & (main_genericstandalone_rtio_core_sed_record6_seqn1[12] != main_genericstandalone_rtio_core_sed_record7_seqn1[12])) ? main_genericstandalone_rtio_core_sed_record6_seqn1[12] : (main_genericstandalone_rtio_core_sed_record6_seqn1 < main_genericstandalone_rtio_core_sed_record7_seqn1))) begin
			main_genericstandalone_rtio_core_sed_record6_rec_valid <= main_genericstandalone_rtio_core_sed_record7_valid0;
			main_genericstandalone_rtio_core_sed_record6_rec_seqn <= main_genericstandalone_rtio_core_sed_record7_seqn1;
			main_genericstandalone_rtio_core_sed_record6_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record7_replace_occured;
			main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record7_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record7_payload_channel1;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record7_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_address <= main_genericstandalone_rtio_core_sed_record7_payload_address1;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_data <= main_genericstandalone_rtio_core_sed_record7_payload_data1;
			main_genericstandalone_rtio_core_sed_record7_rec_valid <= main_genericstandalone_rtio_core_sed_record6_valid0;
			main_genericstandalone_rtio_core_sed_record7_rec_seqn <= main_genericstandalone_rtio_core_sed_record6_seqn1;
			main_genericstandalone_rtio_core_sed_record7_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record6_replace_occured;
			main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record6_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record6_payload_channel1;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record6_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_address <= main_genericstandalone_rtio_core_sed_record6_payload_address1;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_data <= main_genericstandalone_rtio_core_sed_record6_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record6_rec_valid <= main_genericstandalone_rtio_core_sed_record6_valid0;
			main_genericstandalone_rtio_core_sed_record6_rec_seqn <= main_genericstandalone_rtio_core_sed_record6_seqn1;
			main_genericstandalone_rtio_core_sed_record6_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record6_replace_occured;
			main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record6_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record6_payload_channel1;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record6_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_address <= main_genericstandalone_rtio_core_sed_record6_payload_address1;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_data <= main_genericstandalone_rtio_core_sed_record6_payload_data1;
			main_genericstandalone_rtio_core_sed_record7_rec_valid <= main_genericstandalone_rtio_core_sed_record7_valid0;
			main_genericstandalone_rtio_core_sed_record7_rec_seqn <= main_genericstandalone_rtio_core_sed_record7_seqn1;
			main_genericstandalone_rtio_core_sed_record7_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record7_replace_occured;
			main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record7_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record7_payload_channel1;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record7_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_address <= main_genericstandalone_rtio_core_sed_record7_payload_address1;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_data <= main_genericstandalone_rtio_core_sed_record7_payload_data1;
		end
		main_genericstandalone_rtio_core_sed_record6_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference3;
		main_genericstandalone_rtio_core_sed_record7_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record6_valid0), main_genericstandalone_rtio_core_sed_record6_payload_channel1} < {(~main_genericstandalone_rtio_core_sed_record7_valid0), main_genericstandalone_rtio_core_sed_record7_payload_channel1})) begin
			main_genericstandalone_rtio_core_sed_record6_rec_valid <= main_genericstandalone_rtio_core_sed_record6_valid0;
			main_genericstandalone_rtio_core_sed_record6_rec_seqn <= main_genericstandalone_rtio_core_sed_record6_seqn1;
			main_genericstandalone_rtio_core_sed_record6_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record6_replace_occured;
			main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record6_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record6_payload_channel1;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record6_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_address <= main_genericstandalone_rtio_core_sed_record6_payload_address1;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_data <= main_genericstandalone_rtio_core_sed_record6_payload_data1;
			main_genericstandalone_rtio_core_sed_record7_rec_valid <= main_genericstandalone_rtio_core_sed_record7_valid0;
			main_genericstandalone_rtio_core_sed_record7_rec_seqn <= main_genericstandalone_rtio_core_sed_record7_seqn1;
			main_genericstandalone_rtio_core_sed_record7_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record7_replace_occured;
			main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record7_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record7_payload_channel1;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record7_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_address <= main_genericstandalone_rtio_core_sed_record7_payload_address1;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_data <= main_genericstandalone_rtio_core_sed_record7_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record6_rec_valid <= main_genericstandalone_rtio_core_sed_record7_valid0;
			main_genericstandalone_rtio_core_sed_record6_rec_seqn <= main_genericstandalone_rtio_core_sed_record7_seqn1;
			main_genericstandalone_rtio_core_sed_record6_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record7_replace_occured;
			main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record7_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record7_payload_channel1;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record7_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_address <= main_genericstandalone_rtio_core_sed_record7_payload_address1;
			main_genericstandalone_rtio_core_sed_record6_rec_payload_data <= main_genericstandalone_rtio_core_sed_record7_payload_data1;
			main_genericstandalone_rtio_core_sed_record7_rec_valid <= main_genericstandalone_rtio_core_sed_record6_valid0;
			main_genericstandalone_rtio_core_sed_record7_rec_seqn <= main_genericstandalone_rtio_core_sed_record6_seqn1;
			main_genericstandalone_rtio_core_sed_record7_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record6_replace_occured;
			main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record6_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record6_payload_channel1;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record6_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_address <= main_genericstandalone_rtio_core_sed_record6_payload_address1;
			main_genericstandalone_rtio_core_sed_record7_rec_payload_data <= main_genericstandalone_rtio_core_sed_record6_payload_data1;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record8_valid0), main_genericstandalone_rtio_core_sed_record8_payload_channel1} == {(~main_genericstandalone_rtio_core_sed_record9_valid0), main_genericstandalone_rtio_core_sed_record9_payload_channel1})) begin
		if (((((main_genericstandalone_rtio_core_sed_record8_seqn1[11] == main_genericstandalone_rtio_core_sed_record8_seqn1[12]) & (main_genericstandalone_rtio_core_sed_record9_seqn1[11] == main_genericstandalone_rtio_core_sed_record9_seqn1[12])) & (main_genericstandalone_rtio_core_sed_record8_seqn1[12] != main_genericstandalone_rtio_core_sed_record9_seqn1[12])) ? main_genericstandalone_rtio_core_sed_record8_seqn1[12] : (main_genericstandalone_rtio_core_sed_record8_seqn1 < main_genericstandalone_rtio_core_sed_record9_seqn1))) begin
			main_genericstandalone_rtio_core_sed_record8_rec_valid <= main_genericstandalone_rtio_core_sed_record9_valid0;
			main_genericstandalone_rtio_core_sed_record8_rec_seqn <= main_genericstandalone_rtio_core_sed_record9_seqn1;
			main_genericstandalone_rtio_core_sed_record8_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record9_replace_occured;
			main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record9_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record9_payload_channel1;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record9_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_address <= main_genericstandalone_rtio_core_sed_record9_payload_address1;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_data <= main_genericstandalone_rtio_core_sed_record9_payload_data1;
			main_genericstandalone_rtio_core_sed_record9_rec_valid <= main_genericstandalone_rtio_core_sed_record8_valid0;
			main_genericstandalone_rtio_core_sed_record9_rec_seqn <= main_genericstandalone_rtio_core_sed_record8_seqn1;
			main_genericstandalone_rtio_core_sed_record9_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record8_replace_occured;
			main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record8_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record8_payload_channel1;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record8_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_address <= main_genericstandalone_rtio_core_sed_record8_payload_address1;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_data <= main_genericstandalone_rtio_core_sed_record8_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record8_rec_valid <= main_genericstandalone_rtio_core_sed_record8_valid0;
			main_genericstandalone_rtio_core_sed_record8_rec_seqn <= main_genericstandalone_rtio_core_sed_record8_seqn1;
			main_genericstandalone_rtio_core_sed_record8_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record8_replace_occured;
			main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record8_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record8_payload_channel1;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record8_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_address <= main_genericstandalone_rtio_core_sed_record8_payload_address1;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_data <= main_genericstandalone_rtio_core_sed_record8_payload_data1;
			main_genericstandalone_rtio_core_sed_record9_rec_valid <= main_genericstandalone_rtio_core_sed_record9_valid0;
			main_genericstandalone_rtio_core_sed_record9_rec_seqn <= main_genericstandalone_rtio_core_sed_record9_seqn1;
			main_genericstandalone_rtio_core_sed_record9_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record9_replace_occured;
			main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record9_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record9_payload_channel1;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record9_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_address <= main_genericstandalone_rtio_core_sed_record9_payload_address1;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_data <= main_genericstandalone_rtio_core_sed_record9_payload_data1;
		end
		main_genericstandalone_rtio_core_sed_record8_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference4;
		main_genericstandalone_rtio_core_sed_record9_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record8_valid0), main_genericstandalone_rtio_core_sed_record8_payload_channel1} < {(~main_genericstandalone_rtio_core_sed_record9_valid0), main_genericstandalone_rtio_core_sed_record9_payload_channel1})) begin
			main_genericstandalone_rtio_core_sed_record8_rec_valid <= main_genericstandalone_rtio_core_sed_record8_valid0;
			main_genericstandalone_rtio_core_sed_record8_rec_seqn <= main_genericstandalone_rtio_core_sed_record8_seqn1;
			main_genericstandalone_rtio_core_sed_record8_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record8_replace_occured;
			main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record8_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record8_payload_channel1;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record8_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_address <= main_genericstandalone_rtio_core_sed_record8_payload_address1;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_data <= main_genericstandalone_rtio_core_sed_record8_payload_data1;
			main_genericstandalone_rtio_core_sed_record9_rec_valid <= main_genericstandalone_rtio_core_sed_record9_valid0;
			main_genericstandalone_rtio_core_sed_record9_rec_seqn <= main_genericstandalone_rtio_core_sed_record9_seqn1;
			main_genericstandalone_rtio_core_sed_record9_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record9_replace_occured;
			main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record9_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record9_payload_channel1;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record9_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_address <= main_genericstandalone_rtio_core_sed_record9_payload_address1;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_data <= main_genericstandalone_rtio_core_sed_record9_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record8_rec_valid <= main_genericstandalone_rtio_core_sed_record9_valid0;
			main_genericstandalone_rtio_core_sed_record8_rec_seqn <= main_genericstandalone_rtio_core_sed_record9_seqn1;
			main_genericstandalone_rtio_core_sed_record8_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record9_replace_occured;
			main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record9_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record9_payload_channel1;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record9_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_address <= main_genericstandalone_rtio_core_sed_record9_payload_address1;
			main_genericstandalone_rtio_core_sed_record8_rec_payload_data <= main_genericstandalone_rtio_core_sed_record9_payload_data1;
			main_genericstandalone_rtio_core_sed_record9_rec_valid <= main_genericstandalone_rtio_core_sed_record8_valid0;
			main_genericstandalone_rtio_core_sed_record9_rec_seqn <= main_genericstandalone_rtio_core_sed_record8_seqn1;
			main_genericstandalone_rtio_core_sed_record9_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record8_replace_occured;
			main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record8_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record8_payload_channel1;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record8_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_address <= main_genericstandalone_rtio_core_sed_record8_payload_address1;
			main_genericstandalone_rtio_core_sed_record9_rec_payload_data <= main_genericstandalone_rtio_core_sed_record8_payload_data1;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record10_valid0), main_genericstandalone_rtio_core_sed_record10_payload_channel1} == {(~main_genericstandalone_rtio_core_sed_record11_valid0), main_genericstandalone_rtio_core_sed_record11_payload_channel1})) begin
		if (((((main_genericstandalone_rtio_core_sed_record10_seqn1[11] == main_genericstandalone_rtio_core_sed_record10_seqn1[12]) & (main_genericstandalone_rtio_core_sed_record11_seqn1[11] == main_genericstandalone_rtio_core_sed_record11_seqn1[12])) & (main_genericstandalone_rtio_core_sed_record10_seqn1[12] != main_genericstandalone_rtio_core_sed_record11_seqn1[12])) ? main_genericstandalone_rtio_core_sed_record10_seqn1[12] : (main_genericstandalone_rtio_core_sed_record10_seqn1 < main_genericstandalone_rtio_core_sed_record11_seqn1))) begin
			main_genericstandalone_rtio_core_sed_record10_rec_valid <= main_genericstandalone_rtio_core_sed_record11_valid0;
			main_genericstandalone_rtio_core_sed_record10_rec_seqn <= main_genericstandalone_rtio_core_sed_record11_seqn1;
			main_genericstandalone_rtio_core_sed_record10_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record11_replace_occured;
			main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record11_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record11_payload_channel1;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record11_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_address <= main_genericstandalone_rtio_core_sed_record11_payload_address1;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_data <= main_genericstandalone_rtio_core_sed_record11_payload_data1;
			main_genericstandalone_rtio_core_sed_record11_rec_valid <= main_genericstandalone_rtio_core_sed_record10_valid0;
			main_genericstandalone_rtio_core_sed_record11_rec_seqn <= main_genericstandalone_rtio_core_sed_record10_seqn1;
			main_genericstandalone_rtio_core_sed_record11_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record10_replace_occured;
			main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record10_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record10_payload_channel1;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record10_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_address <= main_genericstandalone_rtio_core_sed_record10_payload_address1;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_data <= main_genericstandalone_rtio_core_sed_record10_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record10_rec_valid <= main_genericstandalone_rtio_core_sed_record10_valid0;
			main_genericstandalone_rtio_core_sed_record10_rec_seqn <= main_genericstandalone_rtio_core_sed_record10_seqn1;
			main_genericstandalone_rtio_core_sed_record10_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record10_replace_occured;
			main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record10_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record10_payload_channel1;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record10_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_address <= main_genericstandalone_rtio_core_sed_record10_payload_address1;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_data <= main_genericstandalone_rtio_core_sed_record10_payload_data1;
			main_genericstandalone_rtio_core_sed_record11_rec_valid <= main_genericstandalone_rtio_core_sed_record11_valid0;
			main_genericstandalone_rtio_core_sed_record11_rec_seqn <= main_genericstandalone_rtio_core_sed_record11_seqn1;
			main_genericstandalone_rtio_core_sed_record11_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record11_replace_occured;
			main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record11_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record11_payload_channel1;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record11_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_address <= main_genericstandalone_rtio_core_sed_record11_payload_address1;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_data <= main_genericstandalone_rtio_core_sed_record11_payload_data1;
		end
		main_genericstandalone_rtio_core_sed_record10_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference5;
		main_genericstandalone_rtio_core_sed_record11_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record10_valid0), main_genericstandalone_rtio_core_sed_record10_payload_channel1} < {(~main_genericstandalone_rtio_core_sed_record11_valid0), main_genericstandalone_rtio_core_sed_record11_payload_channel1})) begin
			main_genericstandalone_rtio_core_sed_record10_rec_valid <= main_genericstandalone_rtio_core_sed_record10_valid0;
			main_genericstandalone_rtio_core_sed_record10_rec_seqn <= main_genericstandalone_rtio_core_sed_record10_seqn1;
			main_genericstandalone_rtio_core_sed_record10_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record10_replace_occured;
			main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record10_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record10_payload_channel1;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record10_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_address <= main_genericstandalone_rtio_core_sed_record10_payload_address1;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_data <= main_genericstandalone_rtio_core_sed_record10_payload_data1;
			main_genericstandalone_rtio_core_sed_record11_rec_valid <= main_genericstandalone_rtio_core_sed_record11_valid0;
			main_genericstandalone_rtio_core_sed_record11_rec_seqn <= main_genericstandalone_rtio_core_sed_record11_seqn1;
			main_genericstandalone_rtio_core_sed_record11_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record11_replace_occured;
			main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record11_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record11_payload_channel1;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record11_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_address <= main_genericstandalone_rtio_core_sed_record11_payload_address1;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_data <= main_genericstandalone_rtio_core_sed_record11_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record10_rec_valid <= main_genericstandalone_rtio_core_sed_record11_valid0;
			main_genericstandalone_rtio_core_sed_record10_rec_seqn <= main_genericstandalone_rtio_core_sed_record11_seqn1;
			main_genericstandalone_rtio_core_sed_record10_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record11_replace_occured;
			main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record11_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record11_payload_channel1;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record11_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_address <= main_genericstandalone_rtio_core_sed_record11_payload_address1;
			main_genericstandalone_rtio_core_sed_record10_rec_payload_data <= main_genericstandalone_rtio_core_sed_record11_payload_data1;
			main_genericstandalone_rtio_core_sed_record11_rec_valid <= main_genericstandalone_rtio_core_sed_record10_valid0;
			main_genericstandalone_rtio_core_sed_record11_rec_seqn <= main_genericstandalone_rtio_core_sed_record10_seqn1;
			main_genericstandalone_rtio_core_sed_record11_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record10_replace_occured;
			main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record10_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record10_payload_channel1;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record10_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_address <= main_genericstandalone_rtio_core_sed_record10_payload_address1;
			main_genericstandalone_rtio_core_sed_record11_rec_payload_data <= main_genericstandalone_rtio_core_sed_record10_payload_data1;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record12_valid0), main_genericstandalone_rtio_core_sed_record12_payload_channel1} == {(~main_genericstandalone_rtio_core_sed_record13_valid0), main_genericstandalone_rtio_core_sed_record13_payload_channel1})) begin
		if (((((main_genericstandalone_rtio_core_sed_record12_seqn1[11] == main_genericstandalone_rtio_core_sed_record12_seqn1[12]) & (main_genericstandalone_rtio_core_sed_record13_seqn1[11] == main_genericstandalone_rtio_core_sed_record13_seqn1[12])) & (main_genericstandalone_rtio_core_sed_record12_seqn1[12] != main_genericstandalone_rtio_core_sed_record13_seqn1[12])) ? main_genericstandalone_rtio_core_sed_record12_seqn1[12] : (main_genericstandalone_rtio_core_sed_record12_seqn1 < main_genericstandalone_rtio_core_sed_record13_seqn1))) begin
			main_genericstandalone_rtio_core_sed_record12_rec_valid <= main_genericstandalone_rtio_core_sed_record13_valid0;
			main_genericstandalone_rtio_core_sed_record12_rec_seqn <= main_genericstandalone_rtio_core_sed_record13_seqn1;
			main_genericstandalone_rtio_core_sed_record12_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record13_replace_occured;
			main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record13_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record13_payload_channel1;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record13_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_address <= main_genericstandalone_rtio_core_sed_record13_payload_address1;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_data <= main_genericstandalone_rtio_core_sed_record13_payload_data1;
			main_genericstandalone_rtio_core_sed_record13_rec_valid <= main_genericstandalone_rtio_core_sed_record12_valid0;
			main_genericstandalone_rtio_core_sed_record13_rec_seqn <= main_genericstandalone_rtio_core_sed_record12_seqn1;
			main_genericstandalone_rtio_core_sed_record13_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record12_replace_occured;
			main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record12_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record12_payload_channel1;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record12_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_address <= main_genericstandalone_rtio_core_sed_record12_payload_address1;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_data <= main_genericstandalone_rtio_core_sed_record12_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record12_rec_valid <= main_genericstandalone_rtio_core_sed_record12_valid0;
			main_genericstandalone_rtio_core_sed_record12_rec_seqn <= main_genericstandalone_rtio_core_sed_record12_seqn1;
			main_genericstandalone_rtio_core_sed_record12_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record12_replace_occured;
			main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record12_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record12_payload_channel1;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record12_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_address <= main_genericstandalone_rtio_core_sed_record12_payload_address1;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_data <= main_genericstandalone_rtio_core_sed_record12_payload_data1;
			main_genericstandalone_rtio_core_sed_record13_rec_valid <= main_genericstandalone_rtio_core_sed_record13_valid0;
			main_genericstandalone_rtio_core_sed_record13_rec_seqn <= main_genericstandalone_rtio_core_sed_record13_seqn1;
			main_genericstandalone_rtio_core_sed_record13_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record13_replace_occured;
			main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record13_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record13_payload_channel1;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record13_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_address <= main_genericstandalone_rtio_core_sed_record13_payload_address1;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_data <= main_genericstandalone_rtio_core_sed_record13_payload_data1;
		end
		main_genericstandalone_rtio_core_sed_record12_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference6;
		main_genericstandalone_rtio_core_sed_record13_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record12_valid0), main_genericstandalone_rtio_core_sed_record12_payload_channel1} < {(~main_genericstandalone_rtio_core_sed_record13_valid0), main_genericstandalone_rtio_core_sed_record13_payload_channel1})) begin
			main_genericstandalone_rtio_core_sed_record12_rec_valid <= main_genericstandalone_rtio_core_sed_record12_valid0;
			main_genericstandalone_rtio_core_sed_record12_rec_seqn <= main_genericstandalone_rtio_core_sed_record12_seqn1;
			main_genericstandalone_rtio_core_sed_record12_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record12_replace_occured;
			main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record12_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record12_payload_channel1;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record12_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_address <= main_genericstandalone_rtio_core_sed_record12_payload_address1;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_data <= main_genericstandalone_rtio_core_sed_record12_payload_data1;
			main_genericstandalone_rtio_core_sed_record13_rec_valid <= main_genericstandalone_rtio_core_sed_record13_valid0;
			main_genericstandalone_rtio_core_sed_record13_rec_seqn <= main_genericstandalone_rtio_core_sed_record13_seqn1;
			main_genericstandalone_rtio_core_sed_record13_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record13_replace_occured;
			main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record13_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record13_payload_channel1;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record13_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_address <= main_genericstandalone_rtio_core_sed_record13_payload_address1;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_data <= main_genericstandalone_rtio_core_sed_record13_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record12_rec_valid <= main_genericstandalone_rtio_core_sed_record13_valid0;
			main_genericstandalone_rtio_core_sed_record12_rec_seqn <= main_genericstandalone_rtio_core_sed_record13_seqn1;
			main_genericstandalone_rtio_core_sed_record12_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record13_replace_occured;
			main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record13_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record13_payload_channel1;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record13_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_address <= main_genericstandalone_rtio_core_sed_record13_payload_address1;
			main_genericstandalone_rtio_core_sed_record12_rec_payload_data <= main_genericstandalone_rtio_core_sed_record13_payload_data1;
			main_genericstandalone_rtio_core_sed_record13_rec_valid <= main_genericstandalone_rtio_core_sed_record12_valid0;
			main_genericstandalone_rtio_core_sed_record13_rec_seqn <= main_genericstandalone_rtio_core_sed_record12_seqn1;
			main_genericstandalone_rtio_core_sed_record13_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record12_replace_occured;
			main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record12_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record12_payload_channel1;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record12_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_address <= main_genericstandalone_rtio_core_sed_record12_payload_address1;
			main_genericstandalone_rtio_core_sed_record13_rec_payload_data <= main_genericstandalone_rtio_core_sed_record12_payload_data1;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record14_valid0), main_genericstandalone_rtio_core_sed_record14_payload_channel1} == {(~main_genericstandalone_rtio_core_sed_record15_valid0), main_genericstandalone_rtio_core_sed_record15_payload_channel1})) begin
		if (((((main_genericstandalone_rtio_core_sed_record14_seqn1[11] == main_genericstandalone_rtio_core_sed_record14_seqn1[12]) & (main_genericstandalone_rtio_core_sed_record15_seqn1[11] == main_genericstandalone_rtio_core_sed_record15_seqn1[12])) & (main_genericstandalone_rtio_core_sed_record14_seqn1[12] != main_genericstandalone_rtio_core_sed_record15_seqn1[12])) ? main_genericstandalone_rtio_core_sed_record14_seqn1[12] : (main_genericstandalone_rtio_core_sed_record14_seqn1 < main_genericstandalone_rtio_core_sed_record15_seqn1))) begin
			main_genericstandalone_rtio_core_sed_record14_rec_valid <= main_genericstandalone_rtio_core_sed_record15_valid0;
			main_genericstandalone_rtio_core_sed_record14_rec_seqn <= main_genericstandalone_rtio_core_sed_record15_seqn1;
			main_genericstandalone_rtio_core_sed_record14_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record15_replace_occured;
			main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record15_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record15_payload_channel1;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record15_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_address <= main_genericstandalone_rtio_core_sed_record15_payload_address1;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_data <= main_genericstandalone_rtio_core_sed_record15_payload_data1;
			main_genericstandalone_rtio_core_sed_record15_rec_valid <= main_genericstandalone_rtio_core_sed_record14_valid0;
			main_genericstandalone_rtio_core_sed_record15_rec_seqn <= main_genericstandalone_rtio_core_sed_record14_seqn1;
			main_genericstandalone_rtio_core_sed_record15_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record14_replace_occured;
			main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record14_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record14_payload_channel1;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record14_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_address <= main_genericstandalone_rtio_core_sed_record14_payload_address1;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_data <= main_genericstandalone_rtio_core_sed_record14_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record14_rec_valid <= main_genericstandalone_rtio_core_sed_record14_valid0;
			main_genericstandalone_rtio_core_sed_record14_rec_seqn <= main_genericstandalone_rtio_core_sed_record14_seqn1;
			main_genericstandalone_rtio_core_sed_record14_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record14_replace_occured;
			main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record14_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record14_payload_channel1;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record14_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_address <= main_genericstandalone_rtio_core_sed_record14_payload_address1;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_data <= main_genericstandalone_rtio_core_sed_record14_payload_data1;
			main_genericstandalone_rtio_core_sed_record15_rec_valid <= main_genericstandalone_rtio_core_sed_record15_valid0;
			main_genericstandalone_rtio_core_sed_record15_rec_seqn <= main_genericstandalone_rtio_core_sed_record15_seqn1;
			main_genericstandalone_rtio_core_sed_record15_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record15_replace_occured;
			main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record15_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record15_payload_channel1;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record15_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_address <= main_genericstandalone_rtio_core_sed_record15_payload_address1;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_data <= main_genericstandalone_rtio_core_sed_record15_payload_data1;
		end
		main_genericstandalone_rtio_core_sed_record14_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference7;
		main_genericstandalone_rtio_core_sed_record15_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record14_valid0), main_genericstandalone_rtio_core_sed_record14_payload_channel1} < {(~main_genericstandalone_rtio_core_sed_record15_valid0), main_genericstandalone_rtio_core_sed_record15_payload_channel1})) begin
			main_genericstandalone_rtio_core_sed_record14_rec_valid <= main_genericstandalone_rtio_core_sed_record14_valid0;
			main_genericstandalone_rtio_core_sed_record14_rec_seqn <= main_genericstandalone_rtio_core_sed_record14_seqn1;
			main_genericstandalone_rtio_core_sed_record14_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record14_replace_occured;
			main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record14_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record14_payload_channel1;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record14_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_address <= main_genericstandalone_rtio_core_sed_record14_payload_address1;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_data <= main_genericstandalone_rtio_core_sed_record14_payload_data1;
			main_genericstandalone_rtio_core_sed_record15_rec_valid <= main_genericstandalone_rtio_core_sed_record15_valid0;
			main_genericstandalone_rtio_core_sed_record15_rec_seqn <= main_genericstandalone_rtio_core_sed_record15_seqn1;
			main_genericstandalone_rtio_core_sed_record15_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record15_replace_occured;
			main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record15_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record15_payload_channel1;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record15_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_address <= main_genericstandalone_rtio_core_sed_record15_payload_address1;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_data <= main_genericstandalone_rtio_core_sed_record15_payload_data1;
		end else begin
			main_genericstandalone_rtio_core_sed_record14_rec_valid <= main_genericstandalone_rtio_core_sed_record15_valid0;
			main_genericstandalone_rtio_core_sed_record14_rec_seqn <= main_genericstandalone_rtio_core_sed_record15_seqn1;
			main_genericstandalone_rtio_core_sed_record14_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record15_replace_occured;
			main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record15_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record15_payload_channel1;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record15_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_address <= main_genericstandalone_rtio_core_sed_record15_payload_address1;
			main_genericstandalone_rtio_core_sed_record14_rec_payload_data <= main_genericstandalone_rtio_core_sed_record15_payload_data1;
			main_genericstandalone_rtio_core_sed_record15_rec_valid <= main_genericstandalone_rtio_core_sed_record14_valid0;
			main_genericstandalone_rtio_core_sed_record15_rec_seqn <= main_genericstandalone_rtio_core_sed_record14_seqn1;
			main_genericstandalone_rtio_core_sed_record15_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record14_replace_occured;
			main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record14_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record14_payload_channel1;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record14_payload_fine_ts0;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_address <= main_genericstandalone_rtio_core_sed_record14_payload_address1;
			main_genericstandalone_rtio_core_sed_record15_rec_payload_data <= main_genericstandalone_rtio_core_sed_record14_payload_data1;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record0_rec_valid), main_genericstandalone_rtio_core_sed_record0_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record2_rec_valid), main_genericstandalone_rtio_core_sed_record2_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record0_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record0_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record2_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record2_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record0_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record2_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record0_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record0_rec_seqn < main_genericstandalone_rtio_core_sed_record2_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record16_rec_valid <= main_genericstandalone_rtio_core_sed_record2_rec_valid;
			main_genericstandalone_rtio_core_sed_record16_rec_seqn <= main_genericstandalone_rtio_core_sed_record2_rec_seqn;
			main_genericstandalone_rtio_core_sed_record16_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record2_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record16_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record2_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_address <= main_genericstandalone_rtio_core_sed_record2_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_data <= main_genericstandalone_rtio_core_sed_record2_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record18_rec_valid <= main_genericstandalone_rtio_core_sed_record0_rec_valid;
			main_genericstandalone_rtio_core_sed_record18_rec_seqn <= main_genericstandalone_rtio_core_sed_record0_rec_seqn;
			main_genericstandalone_rtio_core_sed_record18_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record0_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record0_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_address <= main_genericstandalone_rtio_core_sed_record0_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_data <= main_genericstandalone_rtio_core_sed_record0_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record16_rec_valid <= main_genericstandalone_rtio_core_sed_record0_rec_valid;
			main_genericstandalone_rtio_core_sed_record16_rec_seqn <= main_genericstandalone_rtio_core_sed_record0_rec_seqn;
			main_genericstandalone_rtio_core_sed_record16_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record0_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record16_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record0_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_address <= main_genericstandalone_rtio_core_sed_record0_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_data <= main_genericstandalone_rtio_core_sed_record0_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record18_rec_valid <= main_genericstandalone_rtio_core_sed_record2_rec_valid;
			main_genericstandalone_rtio_core_sed_record18_rec_seqn <= main_genericstandalone_rtio_core_sed_record2_rec_seqn;
			main_genericstandalone_rtio_core_sed_record18_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record2_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record2_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_address <= main_genericstandalone_rtio_core_sed_record2_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_data <= main_genericstandalone_rtio_core_sed_record2_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record16_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record16_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference8;
		main_genericstandalone_rtio_core_sed_record18_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record0_rec_valid), main_genericstandalone_rtio_core_sed_record0_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record2_rec_valid), main_genericstandalone_rtio_core_sed_record2_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record16_rec_valid <= main_genericstandalone_rtio_core_sed_record0_rec_valid;
			main_genericstandalone_rtio_core_sed_record16_rec_seqn <= main_genericstandalone_rtio_core_sed_record0_rec_seqn;
			main_genericstandalone_rtio_core_sed_record16_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record0_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record16_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record0_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_address <= main_genericstandalone_rtio_core_sed_record0_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_data <= main_genericstandalone_rtio_core_sed_record0_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record18_rec_valid <= main_genericstandalone_rtio_core_sed_record2_rec_valid;
			main_genericstandalone_rtio_core_sed_record18_rec_seqn <= main_genericstandalone_rtio_core_sed_record2_rec_seqn;
			main_genericstandalone_rtio_core_sed_record18_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record2_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record2_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_address <= main_genericstandalone_rtio_core_sed_record2_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_data <= main_genericstandalone_rtio_core_sed_record2_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record16_rec_valid <= main_genericstandalone_rtio_core_sed_record2_rec_valid;
			main_genericstandalone_rtio_core_sed_record16_rec_seqn <= main_genericstandalone_rtio_core_sed_record2_rec_seqn;
			main_genericstandalone_rtio_core_sed_record16_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record2_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record16_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record2_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record2_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record2_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_address <= main_genericstandalone_rtio_core_sed_record2_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record16_rec_payload_data <= main_genericstandalone_rtio_core_sed_record2_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record18_rec_valid <= main_genericstandalone_rtio_core_sed_record0_rec_valid;
			main_genericstandalone_rtio_core_sed_record18_rec_seqn <= main_genericstandalone_rtio_core_sed_record0_rec_seqn;
			main_genericstandalone_rtio_core_sed_record18_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record0_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record0_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record0_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record0_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_address <= main_genericstandalone_rtio_core_sed_record0_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record18_rec_payload_data <= main_genericstandalone_rtio_core_sed_record0_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record1_rec_valid), main_genericstandalone_rtio_core_sed_record1_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record3_rec_valid), main_genericstandalone_rtio_core_sed_record3_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record1_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record1_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record3_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record3_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record1_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record3_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record1_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record1_rec_seqn < main_genericstandalone_rtio_core_sed_record3_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record17_rec_valid <= main_genericstandalone_rtio_core_sed_record3_rec_valid;
			main_genericstandalone_rtio_core_sed_record17_rec_seqn <= main_genericstandalone_rtio_core_sed_record3_rec_seqn;
			main_genericstandalone_rtio_core_sed_record17_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record3_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record3_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_address <= main_genericstandalone_rtio_core_sed_record3_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_data <= main_genericstandalone_rtio_core_sed_record3_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record19_rec_valid <= main_genericstandalone_rtio_core_sed_record1_rec_valid;
			main_genericstandalone_rtio_core_sed_record19_rec_seqn <= main_genericstandalone_rtio_core_sed_record1_rec_seqn;
			main_genericstandalone_rtio_core_sed_record19_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record1_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record19_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record1_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_address <= main_genericstandalone_rtio_core_sed_record1_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_data <= main_genericstandalone_rtio_core_sed_record1_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record17_rec_valid <= main_genericstandalone_rtio_core_sed_record1_rec_valid;
			main_genericstandalone_rtio_core_sed_record17_rec_seqn <= main_genericstandalone_rtio_core_sed_record1_rec_seqn;
			main_genericstandalone_rtio_core_sed_record17_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record1_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record1_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_address <= main_genericstandalone_rtio_core_sed_record1_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_data <= main_genericstandalone_rtio_core_sed_record1_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record19_rec_valid <= main_genericstandalone_rtio_core_sed_record3_rec_valid;
			main_genericstandalone_rtio_core_sed_record19_rec_seqn <= main_genericstandalone_rtio_core_sed_record3_rec_seqn;
			main_genericstandalone_rtio_core_sed_record19_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record3_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record19_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record3_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_address <= main_genericstandalone_rtio_core_sed_record3_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_data <= main_genericstandalone_rtio_core_sed_record3_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record17_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference9;
		main_genericstandalone_rtio_core_sed_record19_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record1_rec_valid), main_genericstandalone_rtio_core_sed_record1_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record3_rec_valid), main_genericstandalone_rtio_core_sed_record3_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record17_rec_valid <= main_genericstandalone_rtio_core_sed_record1_rec_valid;
			main_genericstandalone_rtio_core_sed_record17_rec_seqn <= main_genericstandalone_rtio_core_sed_record1_rec_seqn;
			main_genericstandalone_rtio_core_sed_record17_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record1_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record1_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_address <= main_genericstandalone_rtio_core_sed_record1_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_data <= main_genericstandalone_rtio_core_sed_record1_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record19_rec_valid <= main_genericstandalone_rtio_core_sed_record3_rec_valid;
			main_genericstandalone_rtio_core_sed_record19_rec_seqn <= main_genericstandalone_rtio_core_sed_record3_rec_seqn;
			main_genericstandalone_rtio_core_sed_record19_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record3_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record19_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record3_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_address <= main_genericstandalone_rtio_core_sed_record3_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_data <= main_genericstandalone_rtio_core_sed_record3_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record17_rec_valid <= main_genericstandalone_rtio_core_sed_record3_rec_valid;
			main_genericstandalone_rtio_core_sed_record17_rec_seqn <= main_genericstandalone_rtio_core_sed_record3_rec_seqn;
			main_genericstandalone_rtio_core_sed_record17_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record3_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record3_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record3_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record3_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_address <= main_genericstandalone_rtio_core_sed_record3_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record17_rec_payload_data <= main_genericstandalone_rtio_core_sed_record3_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record19_rec_valid <= main_genericstandalone_rtio_core_sed_record1_rec_valid;
			main_genericstandalone_rtio_core_sed_record19_rec_seqn <= main_genericstandalone_rtio_core_sed_record1_rec_seqn;
			main_genericstandalone_rtio_core_sed_record19_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record1_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record19_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record1_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record1_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record1_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_address <= main_genericstandalone_rtio_core_sed_record1_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record19_rec_payload_data <= main_genericstandalone_rtio_core_sed_record1_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record4_rec_valid), main_genericstandalone_rtio_core_sed_record4_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record6_rec_valid), main_genericstandalone_rtio_core_sed_record6_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record4_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record4_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record6_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record6_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record4_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record6_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record4_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record4_rec_seqn < main_genericstandalone_rtio_core_sed_record6_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record20_rec_valid <= main_genericstandalone_rtio_core_sed_record6_rec_valid;
			main_genericstandalone_rtio_core_sed_record20_rec_seqn <= main_genericstandalone_rtio_core_sed_record6_rec_seqn;
			main_genericstandalone_rtio_core_sed_record20_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record6_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record20_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record6_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_address <= main_genericstandalone_rtio_core_sed_record6_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_data <= main_genericstandalone_rtio_core_sed_record6_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record22_rec_valid <= main_genericstandalone_rtio_core_sed_record4_rec_valid;
			main_genericstandalone_rtio_core_sed_record22_rec_seqn <= main_genericstandalone_rtio_core_sed_record4_rec_seqn;
			main_genericstandalone_rtio_core_sed_record22_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record4_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record4_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_address <= main_genericstandalone_rtio_core_sed_record4_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_data <= main_genericstandalone_rtio_core_sed_record4_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record20_rec_valid <= main_genericstandalone_rtio_core_sed_record4_rec_valid;
			main_genericstandalone_rtio_core_sed_record20_rec_seqn <= main_genericstandalone_rtio_core_sed_record4_rec_seqn;
			main_genericstandalone_rtio_core_sed_record20_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record4_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record20_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record4_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_address <= main_genericstandalone_rtio_core_sed_record4_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_data <= main_genericstandalone_rtio_core_sed_record4_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record22_rec_valid <= main_genericstandalone_rtio_core_sed_record6_rec_valid;
			main_genericstandalone_rtio_core_sed_record22_rec_seqn <= main_genericstandalone_rtio_core_sed_record6_rec_seqn;
			main_genericstandalone_rtio_core_sed_record22_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record6_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record6_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_address <= main_genericstandalone_rtio_core_sed_record6_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_data <= main_genericstandalone_rtio_core_sed_record6_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record20_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record20_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference10;
		main_genericstandalone_rtio_core_sed_record22_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record4_rec_valid), main_genericstandalone_rtio_core_sed_record4_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record6_rec_valid), main_genericstandalone_rtio_core_sed_record6_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record20_rec_valid <= main_genericstandalone_rtio_core_sed_record4_rec_valid;
			main_genericstandalone_rtio_core_sed_record20_rec_seqn <= main_genericstandalone_rtio_core_sed_record4_rec_seqn;
			main_genericstandalone_rtio_core_sed_record20_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record4_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record20_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record4_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_address <= main_genericstandalone_rtio_core_sed_record4_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_data <= main_genericstandalone_rtio_core_sed_record4_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record22_rec_valid <= main_genericstandalone_rtio_core_sed_record6_rec_valid;
			main_genericstandalone_rtio_core_sed_record22_rec_seqn <= main_genericstandalone_rtio_core_sed_record6_rec_seqn;
			main_genericstandalone_rtio_core_sed_record22_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record6_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record6_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_address <= main_genericstandalone_rtio_core_sed_record6_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_data <= main_genericstandalone_rtio_core_sed_record6_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record20_rec_valid <= main_genericstandalone_rtio_core_sed_record6_rec_valid;
			main_genericstandalone_rtio_core_sed_record20_rec_seqn <= main_genericstandalone_rtio_core_sed_record6_rec_seqn;
			main_genericstandalone_rtio_core_sed_record20_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record6_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record20_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record6_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record6_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record6_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_address <= main_genericstandalone_rtio_core_sed_record6_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record20_rec_payload_data <= main_genericstandalone_rtio_core_sed_record6_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record22_rec_valid <= main_genericstandalone_rtio_core_sed_record4_rec_valid;
			main_genericstandalone_rtio_core_sed_record22_rec_seqn <= main_genericstandalone_rtio_core_sed_record4_rec_seqn;
			main_genericstandalone_rtio_core_sed_record22_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record4_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record4_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record4_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record4_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_address <= main_genericstandalone_rtio_core_sed_record4_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record22_rec_payload_data <= main_genericstandalone_rtio_core_sed_record4_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record5_rec_valid), main_genericstandalone_rtio_core_sed_record5_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record7_rec_valid), main_genericstandalone_rtio_core_sed_record7_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record5_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record5_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record7_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record7_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record5_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record7_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record5_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record5_rec_seqn < main_genericstandalone_rtio_core_sed_record7_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record21_rec_valid <= main_genericstandalone_rtio_core_sed_record7_rec_valid;
			main_genericstandalone_rtio_core_sed_record21_rec_seqn <= main_genericstandalone_rtio_core_sed_record7_rec_seqn;
			main_genericstandalone_rtio_core_sed_record21_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record7_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record7_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_address <= main_genericstandalone_rtio_core_sed_record7_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_data <= main_genericstandalone_rtio_core_sed_record7_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record23_rec_valid <= main_genericstandalone_rtio_core_sed_record5_rec_valid;
			main_genericstandalone_rtio_core_sed_record23_rec_seqn <= main_genericstandalone_rtio_core_sed_record5_rec_seqn;
			main_genericstandalone_rtio_core_sed_record23_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record5_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record23_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record5_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_address <= main_genericstandalone_rtio_core_sed_record5_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_data <= main_genericstandalone_rtio_core_sed_record5_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record21_rec_valid <= main_genericstandalone_rtio_core_sed_record5_rec_valid;
			main_genericstandalone_rtio_core_sed_record21_rec_seqn <= main_genericstandalone_rtio_core_sed_record5_rec_seqn;
			main_genericstandalone_rtio_core_sed_record21_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record5_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record5_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_address <= main_genericstandalone_rtio_core_sed_record5_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_data <= main_genericstandalone_rtio_core_sed_record5_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record23_rec_valid <= main_genericstandalone_rtio_core_sed_record7_rec_valid;
			main_genericstandalone_rtio_core_sed_record23_rec_seqn <= main_genericstandalone_rtio_core_sed_record7_rec_seqn;
			main_genericstandalone_rtio_core_sed_record23_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record7_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record23_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record7_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_address <= main_genericstandalone_rtio_core_sed_record7_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_data <= main_genericstandalone_rtio_core_sed_record7_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record21_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference11;
		main_genericstandalone_rtio_core_sed_record23_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record5_rec_valid), main_genericstandalone_rtio_core_sed_record5_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record7_rec_valid), main_genericstandalone_rtio_core_sed_record7_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record21_rec_valid <= main_genericstandalone_rtio_core_sed_record5_rec_valid;
			main_genericstandalone_rtio_core_sed_record21_rec_seqn <= main_genericstandalone_rtio_core_sed_record5_rec_seqn;
			main_genericstandalone_rtio_core_sed_record21_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record5_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record5_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_address <= main_genericstandalone_rtio_core_sed_record5_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_data <= main_genericstandalone_rtio_core_sed_record5_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record23_rec_valid <= main_genericstandalone_rtio_core_sed_record7_rec_valid;
			main_genericstandalone_rtio_core_sed_record23_rec_seqn <= main_genericstandalone_rtio_core_sed_record7_rec_seqn;
			main_genericstandalone_rtio_core_sed_record23_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record7_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record23_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record7_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_address <= main_genericstandalone_rtio_core_sed_record7_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_data <= main_genericstandalone_rtio_core_sed_record7_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record21_rec_valid <= main_genericstandalone_rtio_core_sed_record7_rec_valid;
			main_genericstandalone_rtio_core_sed_record21_rec_seqn <= main_genericstandalone_rtio_core_sed_record7_rec_seqn;
			main_genericstandalone_rtio_core_sed_record21_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record7_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record7_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record7_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record7_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_address <= main_genericstandalone_rtio_core_sed_record7_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record21_rec_payload_data <= main_genericstandalone_rtio_core_sed_record7_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record23_rec_valid <= main_genericstandalone_rtio_core_sed_record5_rec_valid;
			main_genericstandalone_rtio_core_sed_record23_rec_seqn <= main_genericstandalone_rtio_core_sed_record5_rec_seqn;
			main_genericstandalone_rtio_core_sed_record23_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record5_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record23_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record5_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record5_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record5_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_address <= main_genericstandalone_rtio_core_sed_record5_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record23_rec_payload_data <= main_genericstandalone_rtio_core_sed_record5_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record8_rec_valid), main_genericstandalone_rtio_core_sed_record8_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record10_rec_valid), main_genericstandalone_rtio_core_sed_record10_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record8_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record8_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record10_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record10_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record8_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record10_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record8_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record8_rec_seqn < main_genericstandalone_rtio_core_sed_record10_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record24_rec_valid <= main_genericstandalone_rtio_core_sed_record10_rec_valid;
			main_genericstandalone_rtio_core_sed_record24_rec_seqn <= main_genericstandalone_rtio_core_sed_record10_rec_seqn;
			main_genericstandalone_rtio_core_sed_record24_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record10_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record24_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record10_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_address <= main_genericstandalone_rtio_core_sed_record10_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_data <= main_genericstandalone_rtio_core_sed_record10_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record26_rec_valid <= main_genericstandalone_rtio_core_sed_record8_rec_valid;
			main_genericstandalone_rtio_core_sed_record26_rec_seqn <= main_genericstandalone_rtio_core_sed_record8_rec_seqn;
			main_genericstandalone_rtio_core_sed_record26_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record8_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record8_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_address <= main_genericstandalone_rtio_core_sed_record8_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_data <= main_genericstandalone_rtio_core_sed_record8_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record24_rec_valid <= main_genericstandalone_rtio_core_sed_record8_rec_valid;
			main_genericstandalone_rtio_core_sed_record24_rec_seqn <= main_genericstandalone_rtio_core_sed_record8_rec_seqn;
			main_genericstandalone_rtio_core_sed_record24_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record8_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record24_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record8_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_address <= main_genericstandalone_rtio_core_sed_record8_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_data <= main_genericstandalone_rtio_core_sed_record8_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record26_rec_valid <= main_genericstandalone_rtio_core_sed_record10_rec_valid;
			main_genericstandalone_rtio_core_sed_record26_rec_seqn <= main_genericstandalone_rtio_core_sed_record10_rec_seqn;
			main_genericstandalone_rtio_core_sed_record26_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record10_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record10_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_address <= main_genericstandalone_rtio_core_sed_record10_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_data <= main_genericstandalone_rtio_core_sed_record10_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record24_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record24_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference12;
		main_genericstandalone_rtio_core_sed_record26_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record8_rec_valid), main_genericstandalone_rtio_core_sed_record8_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record10_rec_valid), main_genericstandalone_rtio_core_sed_record10_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record24_rec_valid <= main_genericstandalone_rtio_core_sed_record8_rec_valid;
			main_genericstandalone_rtio_core_sed_record24_rec_seqn <= main_genericstandalone_rtio_core_sed_record8_rec_seqn;
			main_genericstandalone_rtio_core_sed_record24_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record8_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record24_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record8_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_address <= main_genericstandalone_rtio_core_sed_record8_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_data <= main_genericstandalone_rtio_core_sed_record8_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record26_rec_valid <= main_genericstandalone_rtio_core_sed_record10_rec_valid;
			main_genericstandalone_rtio_core_sed_record26_rec_seqn <= main_genericstandalone_rtio_core_sed_record10_rec_seqn;
			main_genericstandalone_rtio_core_sed_record26_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record10_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record10_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_address <= main_genericstandalone_rtio_core_sed_record10_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_data <= main_genericstandalone_rtio_core_sed_record10_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record24_rec_valid <= main_genericstandalone_rtio_core_sed_record10_rec_valid;
			main_genericstandalone_rtio_core_sed_record24_rec_seqn <= main_genericstandalone_rtio_core_sed_record10_rec_seqn;
			main_genericstandalone_rtio_core_sed_record24_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record10_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record24_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record10_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record10_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record10_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_address <= main_genericstandalone_rtio_core_sed_record10_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record24_rec_payload_data <= main_genericstandalone_rtio_core_sed_record10_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record26_rec_valid <= main_genericstandalone_rtio_core_sed_record8_rec_valid;
			main_genericstandalone_rtio_core_sed_record26_rec_seqn <= main_genericstandalone_rtio_core_sed_record8_rec_seqn;
			main_genericstandalone_rtio_core_sed_record26_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record8_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record8_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record8_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record8_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_address <= main_genericstandalone_rtio_core_sed_record8_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record26_rec_payload_data <= main_genericstandalone_rtio_core_sed_record8_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record9_rec_valid), main_genericstandalone_rtio_core_sed_record9_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record11_rec_valid), main_genericstandalone_rtio_core_sed_record11_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record9_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record9_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record11_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record11_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record9_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record11_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record9_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record9_rec_seqn < main_genericstandalone_rtio_core_sed_record11_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record25_rec_valid <= main_genericstandalone_rtio_core_sed_record11_rec_valid;
			main_genericstandalone_rtio_core_sed_record25_rec_seqn <= main_genericstandalone_rtio_core_sed_record11_rec_seqn;
			main_genericstandalone_rtio_core_sed_record25_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record11_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record11_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_address <= main_genericstandalone_rtio_core_sed_record11_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_data <= main_genericstandalone_rtio_core_sed_record11_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record27_rec_valid <= main_genericstandalone_rtio_core_sed_record9_rec_valid;
			main_genericstandalone_rtio_core_sed_record27_rec_seqn <= main_genericstandalone_rtio_core_sed_record9_rec_seqn;
			main_genericstandalone_rtio_core_sed_record27_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record9_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record27_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record9_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_address <= main_genericstandalone_rtio_core_sed_record9_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_data <= main_genericstandalone_rtio_core_sed_record9_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record25_rec_valid <= main_genericstandalone_rtio_core_sed_record9_rec_valid;
			main_genericstandalone_rtio_core_sed_record25_rec_seqn <= main_genericstandalone_rtio_core_sed_record9_rec_seqn;
			main_genericstandalone_rtio_core_sed_record25_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record9_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record9_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_address <= main_genericstandalone_rtio_core_sed_record9_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_data <= main_genericstandalone_rtio_core_sed_record9_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record27_rec_valid <= main_genericstandalone_rtio_core_sed_record11_rec_valid;
			main_genericstandalone_rtio_core_sed_record27_rec_seqn <= main_genericstandalone_rtio_core_sed_record11_rec_seqn;
			main_genericstandalone_rtio_core_sed_record27_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record11_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record27_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record11_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_address <= main_genericstandalone_rtio_core_sed_record11_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_data <= main_genericstandalone_rtio_core_sed_record11_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record25_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference13;
		main_genericstandalone_rtio_core_sed_record27_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record9_rec_valid), main_genericstandalone_rtio_core_sed_record9_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record11_rec_valid), main_genericstandalone_rtio_core_sed_record11_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record25_rec_valid <= main_genericstandalone_rtio_core_sed_record9_rec_valid;
			main_genericstandalone_rtio_core_sed_record25_rec_seqn <= main_genericstandalone_rtio_core_sed_record9_rec_seqn;
			main_genericstandalone_rtio_core_sed_record25_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record9_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record9_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_address <= main_genericstandalone_rtio_core_sed_record9_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_data <= main_genericstandalone_rtio_core_sed_record9_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record27_rec_valid <= main_genericstandalone_rtio_core_sed_record11_rec_valid;
			main_genericstandalone_rtio_core_sed_record27_rec_seqn <= main_genericstandalone_rtio_core_sed_record11_rec_seqn;
			main_genericstandalone_rtio_core_sed_record27_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record11_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record27_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record11_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_address <= main_genericstandalone_rtio_core_sed_record11_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_data <= main_genericstandalone_rtio_core_sed_record11_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record25_rec_valid <= main_genericstandalone_rtio_core_sed_record11_rec_valid;
			main_genericstandalone_rtio_core_sed_record25_rec_seqn <= main_genericstandalone_rtio_core_sed_record11_rec_seqn;
			main_genericstandalone_rtio_core_sed_record25_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record11_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record11_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record11_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record11_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_address <= main_genericstandalone_rtio_core_sed_record11_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record25_rec_payload_data <= main_genericstandalone_rtio_core_sed_record11_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record27_rec_valid <= main_genericstandalone_rtio_core_sed_record9_rec_valid;
			main_genericstandalone_rtio_core_sed_record27_rec_seqn <= main_genericstandalone_rtio_core_sed_record9_rec_seqn;
			main_genericstandalone_rtio_core_sed_record27_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record9_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record27_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record9_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record9_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record9_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_address <= main_genericstandalone_rtio_core_sed_record9_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record27_rec_payload_data <= main_genericstandalone_rtio_core_sed_record9_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record12_rec_valid), main_genericstandalone_rtio_core_sed_record12_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record14_rec_valid), main_genericstandalone_rtio_core_sed_record14_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record12_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record12_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record14_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record14_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record12_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record14_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record12_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record12_rec_seqn < main_genericstandalone_rtio_core_sed_record14_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record28_rec_valid <= main_genericstandalone_rtio_core_sed_record14_rec_valid;
			main_genericstandalone_rtio_core_sed_record28_rec_seqn <= main_genericstandalone_rtio_core_sed_record14_rec_seqn;
			main_genericstandalone_rtio_core_sed_record28_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record14_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record28_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record14_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_address <= main_genericstandalone_rtio_core_sed_record14_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_data <= main_genericstandalone_rtio_core_sed_record14_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record30_rec_valid <= main_genericstandalone_rtio_core_sed_record12_rec_valid;
			main_genericstandalone_rtio_core_sed_record30_rec_seqn <= main_genericstandalone_rtio_core_sed_record12_rec_seqn;
			main_genericstandalone_rtio_core_sed_record30_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record12_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record12_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_address <= main_genericstandalone_rtio_core_sed_record12_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_data <= main_genericstandalone_rtio_core_sed_record12_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record28_rec_valid <= main_genericstandalone_rtio_core_sed_record12_rec_valid;
			main_genericstandalone_rtio_core_sed_record28_rec_seqn <= main_genericstandalone_rtio_core_sed_record12_rec_seqn;
			main_genericstandalone_rtio_core_sed_record28_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record12_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record28_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record12_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_address <= main_genericstandalone_rtio_core_sed_record12_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_data <= main_genericstandalone_rtio_core_sed_record12_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record30_rec_valid <= main_genericstandalone_rtio_core_sed_record14_rec_valid;
			main_genericstandalone_rtio_core_sed_record30_rec_seqn <= main_genericstandalone_rtio_core_sed_record14_rec_seqn;
			main_genericstandalone_rtio_core_sed_record30_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record14_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record14_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_address <= main_genericstandalone_rtio_core_sed_record14_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_data <= main_genericstandalone_rtio_core_sed_record14_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record28_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record28_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference14;
		main_genericstandalone_rtio_core_sed_record30_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record12_rec_valid), main_genericstandalone_rtio_core_sed_record12_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record14_rec_valid), main_genericstandalone_rtio_core_sed_record14_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record28_rec_valid <= main_genericstandalone_rtio_core_sed_record12_rec_valid;
			main_genericstandalone_rtio_core_sed_record28_rec_seqn <= main_genericstandalone_rtio_core_sed_record12_rec_seqn;
			main_genericstandalone_rtio_core_sed_record28_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record12_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record28_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record12_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_address <= main_genericstandalone_rtio_core_sed_record12_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_data <= main_genericstandalone_rtio_core_sed_record12_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record30_rec_valid <= main_genericstandalone_rtio_core_sed_record14_rec_valid;
			main_genericstandalone_rtio_core_sed_record30_rec_seqn <= main_genericstandalone_rtio_core_sed_record14_rec_seqn;
			main_genericstandalone_rtio_core_sed_record30_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record14_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record14_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_address <= main_genericstandalone_rtio_core_sed_record14_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_data <= main_genericstandalone_rtio_core_sed_record14_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record28_rec_valid <= main_genericstandalone_rtio_core_sed_record14_rec_valid;
			main_genericstandalone_rtio_core_sed_record28_rec_seqn <= main_genericstandalone_rtio_core_sed_record14_rec_seqn;
			main_genericstandalone_rtio_core_sed_record28_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record14_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record28_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record14_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record14_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record14_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_address <= main_genericstandalone_rtio_core_sed_record14_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record28_rec_payload_data <= main_genericstandalone_rtio_core_sed_record14_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record30_rec_valid <= main_genericstandalone_rtio_core_sed_record12_rec_valid;
			main_genericstandalone_rtio_core_sed_record30_rec_seqn <= main_genericstandalone_rtio_core_sed_record12_rec_seqn;
			main_genericstandalone_rtio_core_sed_record30_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record12_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record12_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record12_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record12_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_address <= main_genericstandalone_rtio_core_sed_record12_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record30_rec_payload_data <= main_genericstandalone_rtio_core_sed_record12_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record13_rec_valid), main_genericstandalone_rtio_core_sed_record13_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record15_rec_valid), main_genericstandalone_rtio_core_sed_record15_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record13_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record13_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record15_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record15_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record13_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record15_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record13_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record13_rec_seqn < main_genericstandalone_rtio_core_sed_record15_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record29_rec_valid <= main_genericstandalone_rtio_core_sed_record15_rec_valid;
			main_genericstandalone_rtio_core_sed_record29_rec_seqn <= main_genericstandalone_rtio_core_sed_record15_rec_seqn;
			main_genericstandalone_rtio_core_sed_record29_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record15_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record15_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_address <= main_genericstandalone_rtio_core_sed_record15_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_data <= main_genericstandalone_rtio_core_sed_record15_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record31_rec_valid <= main_genericstandalone_rtio_core_sed_record13_rec_valid;
			main_genericstandalone_rtio_core_sed_record31_rec_seqn <= main_genericstandalone_rtio_core_sed_record13_rec_seqn;
			main_genericstandalone_rtio_core_sed_record31_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record13_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record31_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record13_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_address <= main_genericstandalone_rtio_core_sed_record13_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_data <= main_genericstandalone_rtio_core_sed_record13_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record29_rec_valid <= main_genericstandalone_rtio_core_sed_record13_rec_valid;
			main_genericstandalone_rtio_core_sed_record29_rec_seqn <= main_genericstandalone_rtio_core_sed_record13_rec_seqn;
			main_genericstandalone_rtio_core_sed_record29_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record13_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record13_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_address <= main_genericstandalone_rtio_core_sed_record13_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_data <= main_genericstandalone_rtio_core_sed_record13_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record31_rec_valid <= main_genericstandalone_rtio_core_sed_record15_rec_valid;
			main_genericstandalone_rtio_core_sed_record31_rec_seqn <= main_genericstandalone_rtio_core_sed_record15_rec_seqn;
			main_genericstandalone_rtio_core_sed_record31_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record15_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record31_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record15_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_address <= main_genericstandalone_rtio_core_sed_record15_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_data <= main_genericstandalone_rtio_core_sed_record15_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record29_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference15;
		main_genericstandalone_rtio_core_sed_record31_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record13_rec_valid), main_genericstandalone_rtio_core_sed_record13_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record15_rec_valid), main_genericstandalone_rtio_core_sed_record15_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record29_rec_valid <= main_genericstandalone_rtio_core_sed_record13_rec_valid;
			main_genericstandalone_rtio_core_sed_record29_rec_seqn <= main_genericstandalone_rtio_core_sed_record13_rec_seqn;
			main_genericstandalone_rtio_core_sed_record29_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record13_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record13_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_address <= main_genericstandalone_rtio_core_sed_record13_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_data <= main_genericstandalone_rtio_core_sed_record13_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record31_rec_valid <= main_genericstandalone_rtio_core_sed_record15_rec_valid;
			main_genericstandalone_rtio_core_sed_record31_rec_seqn <= main_genericstandalone_rtio_core_sed_record15_rec_seqn;
			main_genericstandalone_rtio_core_sed_record31_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record15_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record31_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record15_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_address <= main_genericstandalone_rtio_core_sed_record15_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_data <= main_genericstandalone_rtio_core_sed_record15_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record29_rec_valid <= main_genericstandalone_rtio_core_sed_record15_rec_valid;
			main_genericstandalone_rtio_core_sed_record29_rec_seqn <= main_genericstandalone_rtio_core_sed_record15_rec_seqn;
			main_genericstandalone_rtio_core_sed_record29_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record15_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record15_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record15_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record15_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_address <= main_genericstandalone_rtio_core_sed_record15_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record29_rec_payload_data <= main_genericstandalone_rtio_core_sed_record15_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record31_rec_valid <= main_genericstandalone_rtio_core_sed_record13_rec_valid;
			main_genericstandalone_rtio_core_sed_record31_rec_seqn <= main_genericstandalone_rtio_core_sed_record13_rec_seqn;
			main_genericstandalone_rtio_core_sed_record31_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record13_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record31_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record13_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record13_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record13_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_address <= main_genericstandalone_rtio_core_sed_record13_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record31_rec_payload_data <= main_genericstandalone_rtio_core_sed_record13_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record17_rec_valid), main_genericstandalone_rtio_core_sed_record17_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record18_rec_valid), main_genericstandalone_rtio_core_sed_record18_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record17_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record17_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record18_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record18_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record17_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record18_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record17_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record17_rec_seqn < main_genericstandalone_rtio_core_sed_record18_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record33_rec_valid <= main_genericstandalone_rtio_core_sed_record18_rec_valid;
			main_genericstandalone_rtio_core_sed_record33_rec_seqn <= main_genericstandalone_rtio_core_sed_record18_rec_seqn;
			main_genericstandalone_rtio_core_sed_record33_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record18_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record18_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_address <= main_genericstandalone_rtio_core_sed_record18_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_data <= main_genericstandalone_rtio_core_sed_record18_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record34_rec_valid <= main_genericstandalone_rtio_core_sed_record17_rec_valid;
			main_genericstandalone_rtio_core_sed_record34_rec_seqn <= main_genericstandalone_rtio_core_sed_record17_rec_seqn;
			main_genericstandalone_rtio_core_sed_record34_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record17_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record17_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_address <= main_genericstandalone_rtio_core_sed_record17_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_data <= main_genericstandalone_rtio_core_sed_record17_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record33_rec_valid <= main_genericstandalone_rtio_core_sed_record17_rec_valid;
			main_genericstandalone_rtio_core_sed_record33_rec_seqn <= main_genericstandalone_rtio_core_sed_record17_rec_seqn;
			main_genericstandalone_rtio_core_sed_record33_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record17_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record17_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_address <= main_genericstandalone_rtio_core_sed_record17_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_data <= main_genericstandalone_rtio_core_sed_record17_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record34_rec_valid <= main_genericstandalone_rtio_core_sed_record18_rec_valid;
			main_genericstandalone_rtio_core_sed_record34_rec_seqn <= main_genericstandalone_rtio_core_sed_record18_rec_seqn;
			main_genericstandalone_rtio_core_sed_record34_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record18_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record18_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_address <= main_genericstandalone_rtio_core_sed_record18_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_data <= main_genericstandalone_rtio_core_sed_record18_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record33_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference16;
		main_genericstandalone_rtio_core_sed_record34_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record17_rec_valid), main_genericstandalone_rtio_core_sed_record17_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record18_rec_valid), main_genericstandalone_rtio_core_sed_record18_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record33_rec_valid <= main_genericstandalone_rtio_core_sed_record17_rec_valid;
			main_genericstandalone_rtio_core_sed_record33_rec_seqn <= main_genericstandalone_rtio_core_sed_record17_rec_seqn;
			main_genericstandalone_rtio_core_sed_record33_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record17_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record17_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_address <= main_genericstandalone_rtio_core_sed_record17_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_data <= main_genericstandalone_rtio_core_sed_record17_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record34_rec_valid <= main_genericstandalone_rtio_core_sed_record18_rec_valid;
			main_genericstandalone_rtio_core_sed_record34_rec_seqn <= main_genericstandalone_rtio_core_sed_record18_rec_seqn;
			main_genericstandalone_rtio_core_sed_record34_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record18_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record18_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_address <= main_genericstandalone_rtio_core_sed_record18_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_data <= main_genericstandalone_rtio_core_sed_record18_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record33_rec_valid <= main_genericstandalone_rtio_core_sed_record18_rec_valid;
			main_genericstandalone_rtio_core_sed_record33_rec_seqn <= main_genericstandalone_rtio_core_sed_record18_rec_seqn;
			main_genericstandalone_rtio_core_sed_record33_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record18_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record18_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record18_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record18_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_address <= main_genericstandalone_rtio_core_sed_record18_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record33_rec_payload_data <= main_genericstandalone_rtio_core_sed_record18_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record34_rec_valid <= main_genericstandalone_rtio_core_sed_record17_rec_valid;
			main_genericstandalone_rtio_core_sed_record34_rec_seqn <= main_genericstandalone_rtio_core_sed_record17_rec_seqn;
			main_genericstandalone_rtio_core_sed_record34_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record17_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record17_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record17_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record17_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_address <= main_genericstandalone_rtio_core_sed_record17_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record34_rec_payload_data <= main_genericstandalone_rtio_core_sed_record17_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record21_rec_valid), main_genericstandalone_rtio_core_sed_record21_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record22_rec_valid), main_genericstandalone_rtio_core_sed_record22_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record21_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record21_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record22_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record22_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record21_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record22_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record21_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record21_rec_seqn < main_genericstandalone_rtio_core_sed_record22_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record37_rec_valid <= main_genericstandalone_rtio_core_sed_record22_rec_valid;
			main_genericstandalone_rtio_core_sed_record37_rec_seqn <= main_genericstandalone_rtio_core_sed_record22_rec_seqn;
			main_genericstandalone_rtio_core_sed_record37_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record22_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record22_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_address <= main_genericstandalone_rtio_core_sed_record22_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_data <= main_genericstandalone_rtio_core_sed_record22_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record38_rec_valid <= main_genericstandalone_rtio_core_sed_record21_rec_valid;
			main_genericstandalone_rtio_core_sed_record38_rec_seqn <= main_genericstandalone_rtio_core_sed_record21_rec_seqn;
			main_genericstandalone_rtio_core_sed_record38_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record21_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record21_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_address <= main_genericstandalone_rtio_core_sed_record21_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_data <= main_genericstandalone_rtio_core_sed_record21_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record37_rec_valid <= main_genericstandalone_rtio_core_sed_record21_rec_valid;
			main_genericstandalone_rtio_core_sed_record37_rec_seqn <= main_genericstandalone_rtio_core_sed_record21_rec_seqn;
			main_genericstandalone_rtio_core_sed_record37_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record21_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record21_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_address <= main_genericstandalone_rtio_core_sed_record21_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_data <= main_genericstandalone_rtio_core_sed_record21_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record38_rec_valid <= main_genericstandalone_rtio_core_sed_record22_rec_valid;
			main_genericstandalone_rtio_core_sed_record38_rec_seqn <= main_genericstandalone_rtio_core_sed_record22_rec_seqn;
			main_genericstandalone_rtio_core_sed_record38_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record22_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record22_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_address <= main_genericstandalone_rtio_core_sed_record22_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_data <= main_genericstandalone_rtio_core_sed_record22_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record37_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference17;
		main_genericstandalone_rtio_core_sed_record38_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record21_rec_valid), main_genericstandalone_rtio_core_sed_record21_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record22_rec_valid), main_genericstandalone_rtio_core_sed_record22_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record37_rec_valid <= main_genericstandalone_rtio_core_sed_record21_rec_valid;
			main_genericstandalone_rtio_core_sed_record37_rec_seqn <= main_genericstandalone_rtio_core_sed_record21_rec_seqn;
			main_genericstandalone_rtio_core_sed_record37_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record21_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record21_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_address <= main_genericstandalone_rtio_core_sed_record21_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_data <= main_genericstandalone_rtio_core_sed_record21_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record38_rec_valid <= main_genericstandalone_rtio_core_sed_record22_rec_valid;
			main_genericstandalone_rtio_core_sed_record38_rec_seqn <= main_genericstandalone_rtio_core_sed_record22_rec_seqn;
			main_genericstandalone_rtio_core_sed_record38_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record22_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record22_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_address <= main_genericstandalone_rtio_core_sed_record22_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_data <= main_genericstandalone_rtio_core_sed_record22_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record37_rec_valid <= main_genericstandalone_rtio_core_sed_record22_rec_valid;
			main_genericstandalone_rtio_core_sed_record37_rec_seqn <= main_genericstandalone_rtio_core_sed_record22_rec_seqn;
			main_genericstandalone_rtio_core_sed_record37_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record22_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record22_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record22_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record22_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_address <= main_genericstandalone_rtio_core_sed_record22_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record37_rec_payload_data <= main_genericstandalone_rtio_core_sed_record22_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record38_rec_valid <= main_genericstandalone_rtio_core_sed_record21_rec_valid;
			main_genericstandalone_rtio_core_sed_record38_rec_seqn <= main_genericstandalone_rtio_core_sed_record21_rec_seqn;
			main_genericstandalone_rtio_core_sed_record38_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record21_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record21_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record21_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record21_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_address <= main_genericstandalone_rtio_core_sed_record21_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record38_rec_payload_data <= main_genericstandalone_rtio_core_sed_record21_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record25_rec_valid), main_genericstandalone_rtio_core_sed_record25_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record26_rec_valid), main_genericstandalone_rtio_core_sed_record26_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record25_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record25_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record26_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record26_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record25_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record26_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record25_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record25_rec_seqn < main_genericstandalone_rtio_core_sed_record26_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record41_rec_valid <= main_genericstandalone_rtio_core_sed_record26_rec_valid;
			main_genericstandalone_rtio_core_sed_record41_rec_seqn <= main_genericstandalone_rtio_core_sed_record26_rec_seqn;
			main_genericstandalone_rtio_core_sed_record41_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record26_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record26_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_address <= main_genericstandalone_rtio_core_sed_record26_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_data <= main_genericstandalone_rtio_core_sed_record26_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record42_rec_valid <= main_genericstandalone_rtio_core_sed_record25_rec_valid;
			main_genericstandalone_rtio_core_sed_record42_rec_seqn <= main_genericstandalone_rtio_core_sed_record25_rec_seqn;
			main_genericstandalone_rtio_core_sed_record42_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record25_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record25_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_address <= main_genericstandalone_rtio_core_sed_record25_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_data <= main_genericstandalone_rtio_core_sed_record25_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record41_rec_valid <= main_genericstandalone_rtio_core_sed_record25_rec_valid;
			main_genericstandalone_rtio_core_sed_record41_rec_seqn <= main_genericstandalone_rtio_core_sed_record25_rec_seqn;
			main_genericstandalone_rtio_core_sed_record41_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record25_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record25_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_address <= main_genericstandalone_rtio_core_sed_record25_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_data <= main_genericstandalone_rtio_core_sed_record25_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record42_rec_valid <= main_genericstandalone_rtio_core_sed_record26_rec_valid;
			main_genericstandalone_rtio_core_sed_record42_rec_seqn <= main_genericstandalone_rtio_core_sed_record26_rec_seqn;
			main_genericstandalone_rtio_core_sed_record42_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record26_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record26_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_address <= main_genericstandalone_rtio_core_sed_record26_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_data <= main_genericstandalone_rtio_core_sed_record26_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record41_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference18;
		main_genericstandalone_rtio_core_sed_record42_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record25_rec_valid), main_genericstandalone_rtio_core_sed_record25_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record26_rec_valid), main_genericstandalone_rtio_core_sed_record26_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record41_rec_valid <= main_genericstandalone_rtio_core_sed_record25_rec_valid;
			main_genericstandalone_rtio_core_sed_record41_rec_seqn <= main_genericstandalone_rtio_core_sed_record25_rec_seqn;
			main_genericstandalone_rtio_core_sed_record41_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record25_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record25_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_address <= main_genericstandalone_rtio_core_sed_record25_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_data <= main_genericstandalone_rtio_core_sed_record25_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record42_rec_valid <= main_genericstandalone_rtio_core_sed_record26_rec_valid;
			main_genericstandalone_rtio_core_sed_record42_rec_seqn <= main_genericstandalone_rtio_core_sed_record26_rec_seqn;
			main_genericstandalone_rtio_core_sed_record42_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record26_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record26_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_address <= main_genericstandalone_rtio_core_sed_record26_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_data <= main_genericstandalone_rtio_core_sed_record26_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record41_rec_valid <= main_genericstandalone_rtio_core_sed_record26_rec_valid;
			main_genericstandalone_rtio_core_sed_record41_rec_seqn <= main_genericstandalone_rtio_core_sed_record26_rec_seqn;
			main_genericstandalone_rtio_core_sed_record41_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record26_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record26_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record26_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record26_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_address <= main_genericstandalone_rtio_core_sed_record26_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record41_rec_payload_data <= main_genericstandalone_rtio_core_sed_record26_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record42_rec_valid <= main_genericstandalone_rtio_core_sed_record25_rec_valid;
			main_genericstandalone_rtio_core_sed_record42_rec_seqn <= main_genericstandalone_rtio_core_sed_record25_rec_seqn;
			main_genericstandalone_rtio_core_sed_record42_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record25_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record25_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record25_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record25_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_address <= main_genericstandalone_rtio_core_sed_record25_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record42_rec_payload_data <= main_genericstandalone_rtio_core_sed_record25_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record29_rec_valid), main_genericstandalone_rtio_core_sed_record29_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record30_rec_valid), main_genericstandalone_rtio_core_sed_record30_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record29_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record29_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record30_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record30_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record29_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record30_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record29_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record29_rec_seqn < main_genericstandalone_rtio_core_sed_record30_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record45_rec_valid <= main_genericstandalone_rtio_core_sed_record30_rec_valid;
			main_genericstandalone_rtio_core_sed_record45_rec_seqn <= main_genericstandalone_rtio_core_sed_record30_rec_seqn;
			main_genericstandalone_rtio_core_sed_record45_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record30_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record30_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_address <= main_genericstandalone_rtio_core_sed_record30_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_data <= main_genericstandalone_rtio_core_sed_record30_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record46_rec_valid <= main_genericstandalone_rtio_core_sed_record29_rec_valid;
			main_genericstandalone_rtio_core_sed_record46_rec_seqn <= main_genericstandalone_rtio_core_sed_record29_rec_seqn;
			main_genericstandalone_rtio_core_sed_record46_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record29_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record29_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_address <= main_genericstandalone_rtio_core_sed_record29_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_data <= main_genericstandalone_rtio_core_sed_record29_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record45_rec_valid <= main_genericstandalone_rtio_core_sed_record29_rec_valid;
			main_genericstandalone_rtio_core_sed_record45_rec_seqn <= main_genericstandalone_rtio_core_sed_record29_rec_seqn;
			main_genericstandalone_rtio_core_sed_record45_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record29_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record29_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_address <= main_genericstandalone_rtio_core_sed_record29_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_data <= main_genericstandalone_rtio_core_sed_record29_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record46_rec_valid <= main_genericstandalone_rtio_core_sed_record30_rec_valid;
			main_genericstandalone_rtio_core_sed_record46_rec_seqn <= main_genericstandalone_rtio_core_sed_record30_rec_seqn;
			main_genericstandalone_rtio_core_sed_record46_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record30_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record30_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_address <= main_genericstandalone_rtio_core_sed_record30_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_data <= main_genericstandalone_rtio_core_sed_record30_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record45_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference19;
		main_genericstandalone_rtio_core_sed_record46_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record29_rec_valid), main_genericstandalone_rtio_core_sed_record29_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record30_rec_valid), main_genericstandalone_rtio_core_sed_record30_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record45_rec_valid <= main_genericstandalone_rtio_core_sed_record29_rec_valid;
			main_genericstandalone_rtio_core_sed_record45_rec_seqn <= main_genericstandalone_rtio_core_sed_record29_rec_seqn;
			main_genericstandalone_rtio_core_sed_record45_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record29_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record29_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_address <= main_genericstandalone_rtio_core_sed_record29_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_data <= main_genericstandalone_rtio_core_sed_record29_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record46_rec_valid <= main_genericstandalone_rtio_core_sed_record30_rec_valid;
			main_genericstandalone_rtio_core_sed_record46_rec_seqn <= main_genericstandalone_rtio_core_sed_record30_rec_seqn;
			main_genericstandalone_rtio_core_sed_record46_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record30_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record30_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_address <= main_genericstandalone_rtio_core_sed_record30_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_data <= main_genericstandalone_rtio_core_sed_record30_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record45_rec_valid <= main_genericstandalone_rtio_core_sed_record30_rec_valid;
			main_genericstandalone_rtio_core_sed_record45_rec_seqn <= main_genericstandalone_rtio_core_sed_record30_rec_seqn;
			main_genericstandalone_rtio_core_sed_record45_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record30_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record30_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record30_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record30_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_address <= main_genericstandalone_rtio_core_sed_record30_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record45_rec_payload_data <= main_genericstandalone_rtio_core_sed_record30_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record46_rec_valid <= main_genericstandalone_rtio_core_sed_record29_rec_valid;
			main_genericstandalone_rtio_core_sed_record46_rec_seqn <= main_genericstandalone_rtio_core_sed_record29_rec_seqn;
			main_genericstandalone_rtio_core_sed_record46_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record29_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record29_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record29_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record29_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_address <= main_genericstandalone_rtio_core_sed_record29_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record46_rec_payload_data <= main_genericstandalone_rtio_core_sed_record29_rec_payload_data;
		end
	end
	main_genericstandalone_rtio_core_sed_record32_rec_valid <= main_genericstandalone_rtio_core_sed_record16_rec_valid;
	main_genericstandalone_rtio_core_sed_record32_rec_seqn <= main_genericstandalone_rtio_core_sed_record16_rec_seqn;
	main_genericstandalone_rtio_core_sed_record32_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record16_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record32_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record16_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record32_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record16_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record32_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record16_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record32_rec_payload_address <= main_genericstandalone_rtio_core_sed_record16_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record32_rec_payload_data <= main_genericstandalone_rtio_core_sed_record16_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record35_rec_valid <= main_genericstandalone_rtio_core_sed_record19_rec_valid;
	main_genericstandalone_rtio_core_sed_record35_rec_seqn <= main_genericstandalone_rtio_core_sed_record19_rec_seqn;
	main_genericstandalone_rtio_core_sed_record35_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record19_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record35_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record19_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record35_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record19_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record35_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record19_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record35_rec_payload_address <= main_genericstandalone_rtio_core_sed_record19_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record35_rec_payload_data <= main_genericstandalone_rtio_core_sed_record19_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record36_rec_valid <= main_genericstandalone_rtio_core_sed_record20_rec_valid;
	main_genericstandalone_rtio_core_sed_record36_rec_seqn <= main_genericstandalone_rtio_core_sed_record20_rec_seqn;
	main_genericstandalone_rtio_core_sed_record36_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record20_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record36_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record20_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record36_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record20_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record36_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record20_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record36_rec_payload_address <= main_genericstandalone_rtio_core_sed_record20_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record36_rec_payload_data <= main_genericstandalone_rtio_core_sed_record20_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record39_rec_valid <= main_genericstandalone_rtio_core_sed_record23_rec_valid;
	main_genericstandalone_rtio_core_sed_record39_rec_seqn <= main_genericstandalone_rtio_core_sed_record23_rec_seqn;
	main_genericstandalone_rtio_core_sed_record39_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record23_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record39_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record23_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record39_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record23_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record39_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record23_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record39_rec_payload_address <= main_genericstandalone_rtio_core_sed_record23_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record39_rec_payload_data <= main_genericstandalone_rtio_core_sed_record23_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record40_rec_valid <= main_genericstandalone_rtio_core_sed_record24_rec_valid;
	main_genericstandalone_rtio_core_sed_record40_rec_seqn <= main_genericstandalone_rtio_core_sed_record24_rec_seqn;
	main_genericstandalone_rtio_core_sed_record40_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record24_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record40_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record24_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record40_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record24_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record40_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record24_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record40_rec_payload_address <= main_genericstandalone_rtio_core_sed_record24_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record40_rec_payload_data <= main_genericstandalone_rtio_core_sed_record24_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record43_rec_valid <= main_genericstandalone_rtio_core_sed_record27_rec_valid;
	main_genericstandalone_rtio_core_sed_record43_rec_seqn <= main_genericstandalone_rtio_core_sed_record27_rec_seqn;
	main_genericstandalone_rtio_core_sed_record43_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record27_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record43_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record27_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record43_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record27_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record43_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record27_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record43_rec_payload_address <= main_genericstandalone_rtio_core_sed_record27_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record43_rec_payload_data <= main_genericstandalone_rtio_core_sed_record27_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record44_rec_valid <= main_genericstandalone_rtio_core_sed_record28_rec_valid;
	main_genericstandalone_rtio_core_sed_record44_rec_seqn <= main_genericstandalone_rtio_core_sed_record28_rec_seqn;
	main_genericstandalone_rtio_core_sed_record44_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record28_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record44_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record28_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record44_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record28_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record44_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record28_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record44_rec_payload_address <= main_genericstandalone_rtio_core_sed_record28_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record44_rec_payload_data <= main_genericstandalone_rtio_core_sed_record28_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record47_rec_valid <= main_genericstandalone_rtio_core_sed_record31_rec_valid;
	main_genericstandalone_rtio_core_sed_record47_rec_seqn <= main_genericstandalone_rtio_core_sed_record31_rec_seqn;
	main_genericstandalone_rtio_core_sed_record47_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record31_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record47_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record31_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record47_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record31_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record47_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record31_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record47_rec_payload_address <= main_genericstandalone_rtio_core_sed_record31_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record47_rec_payload_data <= main_genericstandalone_rtio_core_sed_record31_rec_payload_data;
	if (({(~main_genericstandalone_rtio_core_sed_record32_rec_valid), main_genericstandalone_rtio_core_sed_record32_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record36_rec_valid), main_genericstandalone_rtio_core_sed_record36_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record32_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record32_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record36_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record36_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record32_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record36_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record32_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record32_rec_seqn < main_genericstandalone_rtio_core_sed_record36_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record48_rec_valid <= main_genericstandalone_rtio_core_sed_record36_rec_valid;
			main_genericstandalone_rtio_core_sed_record48_rec_seqn <= main_genericstandalone_rtio_core_sed_record36_rec_seqn;
			main_genericstandalone_rtio_core_sed_record48_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record36_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record48_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record36_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record36_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record36_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_address <= main_genericstandalone_rtio_core_sed_record36_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_data <= main_genericstandalone_rtio_core_sed_record36_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record52_rec_valid <= main_genericstandalone_rtio_core_sed_record32_rec_valid;
			main_genericstandalone_rtio_core_sed_record52_rec_seqn <= main_genericstandalone_rtio_core_sed_record32_rec_seqn;
			main_genericstandalone_rtio_core_sed_record52_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record32_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record32_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record32_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record32_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_address <= main_genericstandalone_rtio_core_sed_record32_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_data <= main_genericstandalone_rtio_core_sed_record32_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record48_rec_valid <= main_genericstandalone_rtio_core_sed_record32_rec_valid;
			main_genericstandalone_rtio_core_sed_record48_rec_seqn <= main_genericstandalone_rtio_core_sed_record32_rec_seqn;
			main_genericstandalone_rtio_core_sed_record48_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record32_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record48_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record32_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record32_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record32_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_address <= main_genericstandalone_rtio_core_sed_record32_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_data <= main_genericstandalone_rtio_core_sed_record32_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record52_rec_valid <= main_genericstandalone_rtio_core_sed_record36_rec_valid;
			main_genericstandalone_rtio_core_sed_record52_rec_seqn <= main_genericstandalone_rtio_core_sed_record36_rec_seqn;
			main_genericstandalone_rtio_core_sed_record52_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record36_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record36_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record36_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record36_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_address <= main_genericstandalone_rtio_core_sed_record36_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_data <= main_genericstandalone_rtio_core_sed_record36_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record48_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record48_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference20;
		main_genericstandalone_rtio_core_sed_record52_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record32_rec_valid), main_genericstandalone_rtio_core_sed_record32_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record36_rec_valid), main_genericstandalone_rtio_core_sed_record36_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record48_rec_valid <= main_genericstandalone_rtio_core_sed_record32_rec_valid;
			main_genericstandalone_rtio_core_sed_record48_rec_seqn <= main_genericstandalone_rtio_core_sed_record32_rec_seqn;
			main_genericstandalone_rtio_core_sed_record48_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record32_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record48_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record32_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record32_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record32_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_address <= main_genericstandalone_rtio_core_sed_record32_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_data <= main_genericstandalone_rtio_core_sed_record32_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record52_rec_valid <= main_genericstandalone_rtio_core_sed_record36_rec_valid;
			main_genericstandalone_rtio_core_sed_record52_rec_seqn <= main_genericstandalone_rtio_core_sed_record36_rec_seqn;
			main_genericstandalone_rtio_core_sed_record52_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record36_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record36_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record36_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record36_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_address <= main_genericstandalone_rtio_core_sed_record36_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_data <= main_genericstandalone_rtio_core_sed_record36_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record48_rec_valid <= main_genericstandalone_rtio_core_sed_record36_rec_valid;
			main_genericstandalone_rtio_core_sed_record48_rec_seqn <= main_genericstandalone_rtio_core_sed_record36_rec_seqn;
			main_genericstandalone_rtio_core_sed_record48_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record36_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record48_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record36_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record36_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record36_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_address <= main_genericstandalone_rtio_core_sed_record36_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record48_rec_payload_data <= main_genericstandalone_rtio_core_sed_record36_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record52_rec_valid <= main_genericstandalone_rtio_core_sed_record32_rec_valid;
			main_genericstandalone_rtio_core_sed_record52_rec_seqn <= main_genericstandalone_rtio_core_sed_record32_rec_seqn;
			main_genericstandalone_rtio_core_sed_record52_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record32_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record32_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record32_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record32_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_address <= main_genericstandalone_rtio_core_sed_record32_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record52_rec_payload_data <= main_genericstandalone_rtio_core_sed_record32_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record33_rec_valid), main_genericstandalone_rtio_core_sed_record33_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record37_rec_valid), main_genericstandalone_rtio_core_sed_record37_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record33_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record33_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record37_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record37_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record33_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record37_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record33_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record33_rec_seqn < main_genericstandalone_rtio_core_sed_record37_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record49_rec_valid <= main_genericstandalone_rtio_core_sed_record37_rec_valid;
			main_genericstandalone_rtio_core_sed_record49_rec_seqn <= main_genericstandalone_rtio_core_sed_record37_rec_seqn;
			main_genericstandalone_rtio_core_sed_record49_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record37_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record49_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record37_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_address <= main_genericstandalone_rtio_core_sed_record37_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_data <= main_genericstandalone_rtio_core_sed_record37_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record53_rec_valid <= main_genericstandalone_rtio_core_sed_record33_rec_valid;
			main_genericstandalone_rtio_core_sed_record53_rec_seqn <= main_genericstandalone_rtio_core_sed_record33_rec_seqn;
			main_genericstandalone_rtio_core_sed_record53_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record33_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record33_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_address <= main_genericstandalone_rtio_core_sed_record33_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_data <= main_genericstandalone_rtio_core_sed_record33_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record49_rec_valid <= main_genericstandalone_rtio_core_sed_record33_rec_valid;
			main_genericstandalone_rtio_core_sed_record49_rec_seqn <= main_genericstandalone_rtio_core_sed_record33_rec_seqn;
			main_genericstandalone_rtio_core_sed_record49_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record33_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record49_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record33_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_address <= main_genericstandalone_rtio_core_sed_record33_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_data <= main_genericstandalone_rtio_core_sed_record33_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record53_rec_valid <= main_genericstandalone_rtio_core_sed_record37_rec_valid;
			main_genericstandalone_rtio_core_sed_record53_rec_seqn <= main_genericstandalone_rtio_core_sed_record37_rec_seqn;
			main_genericstandalone_rtio_core_sed_record53_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record37_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record37_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_address <= main_genericstandalone_rtio_core_sed_record37_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_data <= main_genericstandalone_rtio_core_sed_record37_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record49_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record49_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference21;
		main_genericstandalone_rtio_core_sed_record53_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record33_rec_valid), main_genericstandalone_rtio_core_sed_record33_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record37_rec_valid), main_genericstandalone_rtio_core_sed_record37_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record49_rec_valid <= main_genericstandalone_rtio_core_sed_record33_rec_valid;
			main_genericstandalone_rtio_core_sed_record49_rec_seqn <= main_genericstandalone_rtio_core_sed_record33_rec_seqn;
			main_genericstandalone_rtio_core_sed_record49_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record33_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record49_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record33_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_address <= main_genericstandalone_rtio_core_sed_record33_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_data <= main_genericstandalone_rtio_core_sed_record33_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record53_rec_valid <= main_genericstandalone_rtio_core_sed_record37_rec_valid;
			main_genericstandalone_rtio_core_sed_record53_rec_seqn <= main_genericstandalone_rtio_core_sed_record37_rec_seqn;
			main_genericstandalone_rtio_core_sed_record53_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record37_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record37_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_address <= main_genericstandalone_rtio_core_sed_record37_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_data <= main_genericstandalone_rtio_core_sed_record37_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record49_rec_valid <= main_genericstandalone_rtio_core_sed_record37_rec_valid;
			main_genericstandalone_rtio_core_sed_record49_rec_seqn <= main_genericstandalone_rtio_core_sed_record37_rec_seqn;
			main_genericstandalone_rtio_core_sed_record49_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record37_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record49_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record37_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record37_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record37_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_address <= main_genericstandalone_rtio_core_sed_record37_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record49_rec_payload_data <= main_genericstandalone_rtio_core_sed_record37_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record53_rec_valid <= main_genericstandalone_rtio_core_sed_record33_rec_valid;
			main_genericstandalone_rtio_core_sed_record53_rec_seqn <= main_genericstandalone_rtio_core_sed_record33_rec_seqn;
			main_genericstandalone_rtio_core_sed_record53_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record33_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record33_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record33_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record33_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_address <= main_genericstandalone_rtio_core_sed_record33_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record53_rec_payload_data <= main_genericstandalone_rtio_core_sed_record33_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record34_rec_valid), main_genericstandalone_rtio_core_sed_record34_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record38_rec_valid), main_genericstandalone_rtio_core_sed_record38_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record34_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record34_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record38_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record38_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record34_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record38_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record34_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record34_rec_seqn < main_genericstandalone_rtio_core_sed_record38_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record50_rec_valid <= main_genericstandalone_rtio_core_sed_record38_rec_valid;
			main_genericstandalone_rtio_core_sed_record50_rec_seqn <= main_genericstandalone_rtio_core_sed_record38_rec_seqn;
			main_genericstandalone_rtio_core_sed_record50_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record38_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record38_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_address <= main_genericstandalone_rtio_core_sed_record38_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_data <= main_genericstandalone_rtio_core_sed_record38_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record54_rec_valid <= main_genericstandalone_rtio_core_sed_record34_rec_valid;
			main_genericstandalone_rtio_core_sed_record54_rec_seqn <= main_genericstandalone_rtio_core_sed_record34_rec_seqn;
			main_genericstandalone_rtio_core_sed_record54_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record34_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record54_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record34_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_address <= main_genericstandalone_rtio_core_sed_record34_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_data <= main_genericstandalone_rtio_core_sed_record34_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record50_rec_valid <= main_genericstandalone_rtio_core_sed_record34_rec_valid;
			main_genericstandalone_rtio_core_sed_record50_rec_seqn <= main_genericstandalone_rtio_core_sed_record34_rec_seqn;
			main_genericstandalone_rtio_core_sed_record50_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record34_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record34_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_address <= main_genericstandalone_rtio_core_sed_record34_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_data <= main_genericstandalone_rtio_core_sed_record34_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record54_rec_valid <= main_genericstandalone_rtio_core_sed_record38_rec_valid;
			main_genericstandalone_rtio_core_sed_record54_rec_seqn <= main_genericstandalone_rtio_core_sed_record38_rec_seqn;
			main_genericstandalone_rtio_core_sed_record54_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record38_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record54_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record38_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_address <= main_genericstandalone_rtio_core_sed_record38_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_data <= main_genericstandalone_rtio_core_sed_record38_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record50_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference22;
		main_genericstandalone_rtio_core_sed_record54_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record34_rec_valid), main_genericstandalone_rtio_core_sed_record34_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record38_rec_valid), main_genericstandalone_rtio_core_sed_record38_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record50_rec_valid <= main_genericstandalone_rtio_core_sed_record34_rec_valid;
			main_genericstandalone_rtio_core_sed_record50_rec_seqn <= main_genericstandalone_rtio_core_sed_record34_rec_seqn;
			main_genericstandalone_rtio_core_sed_record50_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record34_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record34_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_address <= main_genericstandalone_rtio_core_sed_record34_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_data <= main_genericstandalone_rtio_core_sed_record34_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record54_rec_valid <= main_genericstandalone_rtio_core_sed_record38_rec_valid;
			main_genericstandalone_rtio_core_sed_record54_rec_seqn <= main_genericstandalone_rtio_core_sed_record38_rec_seqn;
			main_genericstandalone_rtio_core_sed_record54_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record38_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record54_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record38_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_address <= main_genericstandalone_rtio_core_sed_record38_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_data <= main_genericstandalone_rtio_core_sed_record38_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record50_rec_valid <= main_genericstandalone_rtio_core_sed_record38_rec_valid;
			main_genericstandalone_rtio_core_sed_record50_rec_seqn <= main_genericstandalone_rtio_core_sed_record38_rec_seqn;
			main_genericstandalone_rtio_core_sed_record50_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record38_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record38_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record38_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record38_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_address <= main_genericstandalone_rtio_core_sed_record38_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record50_rec_payload_data <= main_genericstandalone_rtio_core_sed_record38_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record54_rec_valid <= main_genericstandalone_rtio_core_sed_record34_rec_valid;
			main_genericstandalone_rtio_core_sed_record54_rec_seqn <= main_genericstandalone_rtio_core_sed_record34_rec_seqn;
			main_genericstandalone_rtio_core_sed_record54_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record34_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record54_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record34_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record34_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record34_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_address <= main_genericstandalone_rtio_core_sed_record34_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record54_rec_payload_data <= main_genericstandalone_rtio_core_sed_record34_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record35_rec_valid), main_genericstandalone_rtio_core_sed_record35_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record39_rec_valid), main_genericstandalone_rtio_core_sed_record39_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record35_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record35_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record39_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record39_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record35_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record39_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record35_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record35_rec_seqn < main_genericstandalone_rtio_core_sed_record39_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record51_rec_valid <= main_genericstandalone_rtio_core_sed_record39_rec_valid;
			main_genericstandalone_rtio_core_sed_record51_rec_seqn <= main_genericstandalone_rtio_core_sed_record39_rec_seqn;
			main_genericstandalone_rtio_core_sed_record51_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record39_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record39_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record39_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record39_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_address <= main_genericstandalone_rtio_core_sed_record39_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_data <= main_genericstandalone_rtio_core_sed_record39_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record55_rec_valid <= main_genericstandalone_rtio_core_sed_record35_rec_valid;
			main_genericstandalone_rtio_core_sed_record55_rec_seqn <= main_genericstandalone_rtio_core_sed_record35_rec_seqn;
			main_genericstandalone_rtio_core_sed_record55_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record35_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record55_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record35_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record35_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record35_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_address <= main_genericstandalone_rtio_core_sed_record35_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_data <= main_genericstandalone_rtio_core_sed_record35_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record51_rec_valid <= main_genericstandalone_rtio_core_sed_record35_rec_valid;
			main_genericstandalone_rtio_core_sed_record51_rec_seqn <= main_genericstandalone_rtio_core_sed_record35_rec_seqn;
			main_genericstandalone_rtio_core_sed_record51_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record35_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record35_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record35_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record35_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_address <= main_genericstandalone_rtio_core_sed_record35_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_data <= main_genericstandalone_rtio_core_sed_record35_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record55_rec_valid <= main_genericstandalone_rtio_core_sed_record39_rec_valid;
			main_genericstandalone_rtio_core_sed_record55_rec_seqn <= main_genericstandalone_rtio_core_sed_record39_rec_seqn;
			main_genericstandalone_rtio_core_sed_record55_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record39_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record55_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record39_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record39_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record39_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_address <= main_genericstandalone_rtio_core_sed_record39_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_data <= main_genericstandalone_rtio_core_sed_record39_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record51_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference23;
		main_genericstandalone_rtio_core_sed_record55_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record35_rec_valid), main_genericstandalone_rtio_core_sed_record35_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record39_rec_valid), main_genericstandalone_rtio_core_sed_record39_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record51_rec_valid <= main_genericstandalone_rtio_core_sed_record35_rec_valid;
			main_genericstandalone_rtio_core_sed_record51_rec_seqn <= main_genericstandalone_rtio_core_sed_record35_rec_seqn;
			main_genericstandalone_rtio_core_sed_record51_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record35_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record35_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record35_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record35_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_address <= main_genericstandalone_rtio_core_sed_record35_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_data <= main_genericstandalone_rtio_core_sed_record35_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record55_rec_valid <= main_genericstandalone_rtio_core_sed_record39_rec_valid;
			main_genericstandalone_rtio_core_sed_record55_rec_seqn <= main_genericstandalone_rtio_core_sed_record39_rec_seqn;
			main_genericstandalone_rtio_core_sed_record55_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record39_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record55_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record39_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record39_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record39_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_address <= main_genericstandalone_rtio_core_sed_record39_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_data <= main_genericstandalone_rtio_core_sed_record39_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record51_rec_valid <= main_genericstandalone_rtio_core_sed_record39_rec_valid;
			main_genericstandalone_rtio_core_sed_record51_rec_seqn <= main_genericstandalone_rtio_core_sed_record39_rec_seqn;
			main_genericstandalone_rtio_core_sed_record51_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record39_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record39_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record39_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record39_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_address <= main_genericstandalone_rtio_core_sed_record39_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record51_rec_payload_data <= main_genericstandalone_rtio_core_sed_record39_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record55_rec_valid <= main_genericstandalone_rtio_core_sed_record35_rec_valid;
			main_genericstandalone_rtio_core_sed_record55_rec_seqn <= main_genericstandalone_rtio_core_sed_record35_rec_seqn;
			main_genericstandalone_rtio_core_sed_record55_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record35_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record55_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record35_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record35_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record35_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_address <= main_genericstandalone_rtio_core_sed_record35_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record55_rec_payload_data <= main_genericstandalone_rtio_core_sed_record35_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record40_rec_valid), main_genericstandalone_rtio_core_sed_record40_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record44_rec_valid), main_genericstandalone_rtio_core_sed_record44_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record40_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record40_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record44_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record44_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record40_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record44_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record40_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record40_rec_seqn < main_genericstandalone_rtio_core_sed_record44_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record56_rec_valid <= main_genericstandalone_rtio_core_sed_record44_rec_valid;
			main_genericstandalone_rtio_core_sed_record56_rec_seqn <= main_genericstandalone_rtio_core_sed_record44_rec_seqn;
			main_genericstandalone_rtio_core_sed_record56_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record44_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record56_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record44_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record44_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record44_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_address <= main_genericstandalone_rtio_core_sed_record44_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_data <= main_genericstandalone_rtio_core_sed_record44_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record60_rec_valid <= main_genericstandalone_rtio_core_sed_record40_rec_valid;
			main_genericstandalone_rtio_core_sed_record60_rec_seqn <= main_genericstandalone_rtio_core_sed_record40_rec_seqn;
			main_genericstandalone_rtio_core_sed_record60_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record40_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record40_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record40_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record40_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_address <= main_genericstandalone_rtio_core_sed_record40_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_data <= main_genericstandalone_rtio_core_sed_record40_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record56_rec_valid <= main_genericstandalone_rtio_core_sed_record40_rec_valid;
			main_genericstandalone_rtio_core_sed_record56_rec_seqn <= main_genericstandalone_rtio_core_sed_record40_rec_seqn;
			main_genericstandalone_rtio_core_sed_record56_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record40_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record56_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record40_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record40_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record40_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_address <= main_genericstandalone_rtio_core_sed_record40_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_data <= main_genericstandalone_rtio_core_sed_record40_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record60_rec_valid <= main_genericstandalone_rtio_core_sed_record44_rec_valid;
			main_genericstandalone_rtio_core_sed_record60_rec_seqn <= main_genericstandalone_rtio_core_sed_record44_rec_seqn;
			main_genericstandalone_rtio_core_sed_record60_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record44_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record44_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record44_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record44_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_address <= main_genericstandalone_rtio_core_sed_record44_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_data <= main_genericstandalone_rtio_core_sed_record44_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record56_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record56_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference24;
		main_genericstandalone_rtio_core_sed_record60_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record40_rec_valid), main_genericstandalone_rtio_core_sed_record40_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record44_rec_valid), main_genericstandalone_rtio_core_sed_record44_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record56_rec_valid <= main_genericstandalone_rtio_core_sed_record40_rec_valid;
			main_genericstandalone_rtio_core_sed_record56_rec_seqn <= main_genericstandalone_rtio_core_sed_record40_rec_seqn;
			main_genericstandalone_rtio_core_sed_record56_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record40_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record56_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record40_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record40_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record40_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_address <= main_genericstandalone_rtio_core_sed_record40_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_data <= main_genericstandalone_rtio_core_sed_record40_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record60_rec_valid <= main_genericstandalone_rtio_core_sed_record44_rec_valid;
			main_genericstandalone_rtio_core_sed_record60_rec_seqn <= main_genericstandalone_rtio_core_sed_record44_rec_seqn;
			main_genericstandalone_rtio_core_sed_record60_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record44_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record44_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record44_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record44_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_address <= main_genericstandalone_rtio_core_sed_record44_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_data <= main_genericstandalone_rtio_core_sed_record44_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record56_rec_valid <= main_genericstandalone_rtio_core_sed_record44_rec_valid;
			main_genericstandalone_rtio_core_sed_record56_rec_seqn <= main_genericstandalone_rtio_core_sed_record44_rec_seqn;
			main_genericstandalone_rtio_core_sed_record56_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record44_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record56_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record44_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record44_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record44_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_address <= main_genericstandalone_rtio_core_sed_record44_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record56_rec_payload_data <= main_genericstandalone_rtio_core_sed_record44_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record60_rec_valid <= main_genericstandalone_rtio_core_sed_record40_rec_valid;
			main_genericstandalone_rtio_core_sed_record60_rec_seqn <= main_genericstandalone_rtio_core_sed_record40_rec_seqn;
			main_genericstandalone_rtio_core_sed_record60_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record40_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record40_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record40_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record40_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_address <= main_genericstandalone_rtio_core_sed_record40_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record60_rec_payload_data <= main_genericstandalone_rtio_core_sed_record40_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record41_rec_valid), main_genericstandalone_rtio_core_sed_record41_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record45_rec_valid), main_genericstandalone_rtio_core_sed_record45_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record41_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record41_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record45_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record45_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record41_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record45_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record41_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record41_rec_seqn < main_genericstandalone_rtio_core_sed_record45_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record57_rec_valid <= main_genericstandalone_rtio_core_sed_record45_rec_valid;
			main_genericstandalone_rtio_core_sed_record57_rec_seqn <= main_genericstandalone_rtio_core_sed_record45_rec_seqn;
			main_genericstandalone_rtio_core_sed_record57_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record45_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record57_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record45_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_address <= main_genericstandalone_rtio_core_sed_record45_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_data <= main_genericstandalone_rtio_core_sed_record45_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record61_rec_valid <= main_genericstandalone_rtio_core_sed_record41_rec_valid;
			main_genericstandalone_rtio_core_sed_record61_rec_seqn <= main_genericstandalone_rtio_core_sed_record41_rec_seqn;
			main_genericstandalone_rtio_core_sed_record61_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record41_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record41_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_address <= main_genericstandalone_rtio_core_sed_record41_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_data <= main_genericstandalone_rtio_core_sed_record41_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record57_rec_valid <= main_genericstandalone_rtio_core_sed_record41_rec_valid;
			main_genericstandalone_rtio_core_sed_record57_rec_seqn <= main_genericstandalone_rtio_core_sed_record41_rec_seqn;
			main_genericstandalone_rtio_core_sed_record57_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record41_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record57_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record41_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_address <= main_genericstandalone_rtio_core_sed_record41_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_data <= main_genericstandalone_rtio_core_sed_record41_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record61_rec_valid <= main_genericstandalone_rtio_core_sed_record45_rec_valid;
			main_genericstandalone_rtio_core_sed_record61_rec_seqn <= main_genericstandalone_rtio_core_sed_record45_rec_seqn;
			main_genericstandalone_rtio_core_sed_record61_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record45_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record45_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_address <= main_genericstandalone_rtio_core_sed_record45_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_data <= main_genericstandalone_rtio_core_sed_record45_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record57_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record57_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference25;
		main_genericstandalone_rtio_core_sed_record61_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record41_rec_valid), main_genericstandalone_rtio_core_sed_record41_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record45_rec_valid), main_genericstandalone_rtio_core_sed_record45_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record57_rec_valid <= main_genericstandalone_rtio_core_sed_record41_rec_valid;
			main_genericstandalone_rtio_core_sed_record57_rec_seqn <= main_genericstandalone_rtio_core_sed_record41_rec_seqn;
			main_genericstandalone_rtio_core_sed_record57_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record41_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record57_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record41_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_address <= main_genericstandalone_rtio_core_sed_record41_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_data <= main_genericstandalone_rtio_core_sed_record41_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record61_rec_valid <= main_genericstandalone_rtio_core_sed_record45_rec_valid;
			main_genericstandalone_rtio_core_sed_record61_rec_seqn <= main_genericstandalone_rtio_core_sed_record45_rec_seqn;
			main_genericstandalone_rtio_core_sed_record61_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record45_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record45_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_address <= main_genericstandalone_rtio_core_sed_record45_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_data <= main_genericstandalone_rtio_core_sed_record45_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record57_rec_valid <= main_genericstandalone_rtio_core_sed_record45_rec_valid;
			main_genericstandalone_rtio_core_sed_record57_rec_seqn <= main_genericstandalone_rtio_core_sed_record45_rec_seqn;
			main_genericstandalone_rtio_core_sed_record57_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record45_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record57_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record45_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record45_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record45_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_address <= main_genericstandalone_rtio_core_sed_record45_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record57_rec_payload_data <= main_genericstandalone_rtio_core_sed_record45_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record61_rec_valid <= main_genericstandalone_rtio_core_sed_record41_rec_valid;
			main_genericstandalone_rtio_core_sed_record61_rec_seqn <= main_genericstandalone_rtio_core_sed_record41_rec_seqn;
			main_genericstandalone_rtio_core_sed_record61_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record41_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record41_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record41_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record41_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_address <= main_genericstandalone_rtio_core_sed_record41_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record61_rec_payload_data <= main_genericstandalone_rtio_core_sed_record41_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record42_rec_valid), main_genericstandalone_rtio_core_sed_record42_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record46_rec_valid), main_genericstandalone_rtio_core_sed_record46_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record42_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record42_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record46_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record46_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record42_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record46_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record42_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record42_rec_seqn < main_genericstandalone_rtio_core_sed_record46_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record58_rec_valid <= main_genericstandalone_rtio_core_sed_record46_rec_valid;
			main_genericstandalone_rtio_core_sed_record58_rec_seqn <= main_genericstandalone_rtio_core_sed_record46_rec_seqn;
			main_genericstandalone_rtio_core_sed_record58_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record46_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record46_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_address <= main_genericstandalone_rtio_core_sed_record46_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_data <= main_genericstandalone_rtio_core_sed_record46_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record62_rec_valid <= main_genericstandalone_rtio_core_sed_record42_rec_valid;
			main_genericstandalone_rtio_core_sed_record62_rec_seqn <= main_genericstandalone_rtio_core_sed_record42_rec_seqn;
			main_genericstandalone_rtio_core_sed_record62_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record42_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record62_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record42_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_address <= main_genericstandalone_rtio_core_sed_record42_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_data <= main_genericstandalone_rtio_core_sed_record42_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record58_rec_valid <= main_genericstandalone_rtio_core_sed_record42_rec_valid;
			main_genericstandalone_rtio_core_sed_record58_rec_seqn <= main_genericstandalone_rtio_core_sed_record42_rec_seqn;
			main_genericstandalone_rtio_core_sed_record58_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record42_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record42_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_address <= main_genericstandalone_rtio_core_sed_record42_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_data <= main_genericstandalone_rtio_core_sed_record42_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record62_rec_valid <= main_genericstandalone_rtio_core_sed_record46_rec_valid;
			main_genericstandalone_rtio_core_sed_record62_rec_seqn <= main_genericstandalone_rtio_core_sed_record46_rec_seqn;
			main_genericstandalone_rtio_core_sed_record62_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record46_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record62_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record46_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_address <= main_genericstandalone_rtio_core_sed_record46_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_data <= main_genericstandalone_rtio_core_sed_record46_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record58_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference26;
		main_genericstandalone_rtio_core_sed_record62_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record42_rec_valid), main_genericstandalone_rtio_core_sed_record42_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record46_rec_valid), main_genericstandalone_rtio_core_sed_record46_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record58_rec_valid <= main_genericstandalone_rtio_core_sed_record42_rec_valid;
			main_genericstandalone_rtio_core_sed_record58_rec_seqn <= main_genericstandalone_rtio_core_sed_record42_rec_seqn;
			main_genericstandalone_rtio_core_sed_record58_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record42_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record42_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_address <= main_genericstandalone_rtio_core_sed_record42_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_data <= main_genericstandalone_rtio_core_sed_record42_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record62_rec_valid <= main_genericstandalone_rtio_core_sed_record46_rec_valid;
			main_genericstandalone_rtio_core_sed_record62_rec_seqn <= main_genericstandalone_rtio_core_sed_record46_rec_seqn;
			main_genericstandalone_rtio_core_sed_record62_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record46_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record62_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record46_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_address <= main_genericstandalone_rtio_core_sed_record46_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_data <= main_genericstandalone_rtio_core_sed_record46_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record58_rec_valid <= main_genericstandalone_rtio_core_sed_record46_rec_valid;
			main_genericstandalone_rtio_core_sed_record58_rec_seqn <= main_genericstandalone_rtio_core_sed_record46_rec_seqn;
			main_genericstandalone_rtio_core_sed_record58_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record46_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record46_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record46_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record46_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_address <= main_genericstandalone_rtio_core_sed_record46_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record58_rec_payload_data <= main_genericstandalone_rtio_core_sed_record46_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record62_rec_valid <= main_genericstandalone_rtio_core_sed_record42_rec_valid;
			main_genericstandalone_rtio_core_sed_record62_rec_seqn <= main_genericstandalone_rtio_core_sed_record42_rec_seqn;
			main_genericstandalone_rtio_core_sed_record62_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record42_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record62_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record42_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record42_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record42_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_address <= main_genericstandalone_rtio_core_sed_record42_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record62_rec_payload_data <= main_genericstandalone_rtio_core_sed_record42_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record43_rec_valid), main_genericstandalone_rtio_core_sed_record43_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record47_rec_valid), main_genericstandalone_rtio_core_sed_record47_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record43_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record43_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record47_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record47_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record43_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record47_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record43_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record43_rec_seqn < main_genericstandalone_rtio_core_sed_record47_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record59_rec_valid <= main_genericstandalone_rtio_core_sed_record47_rec_valid;
			main_genericstandalone_rtio_core_sed_record59_rec_seqn <= main_genericstandalone_rtio_core_sed_record47_rec_seqn;
			main_genericstandalone_rtio_core_sed_record59_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record47_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record47_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record47_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record47_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_address <= main_genericstandalone_rtio_core_sed_record47_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_data <= main_genericstandalone_rtio_core_sed_record47_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record63_rec_valid <= main_genericstandalone_rtio_core_sed_record43_rec_valid;
			main_genericstandalone_rtio_core_sed_record63_rec_seqn <= main_genericstandalone_rtio_core_sed_record43_rec_seqn;
			main_genericstandalone_rtio_core_sed_record63_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record43_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record63_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record43_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record43_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record43_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_address <= main_genericstandalone_rtio_core_sed_record43_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_data <= main_genericstandalone_rtio_core_sed_record43_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record59_rec_valid <= main_genericstandalone_rtio_core_sed_record43_rec_valid;
			main_genericstandalone_rtio_core_sed_record59_rec_seqn <= main_genericstandalone_rtio_core_sed_record43_rec_seqn;
			main_genericstandalone_rtio_core_sed_record59_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record43_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record43_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record43_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record43_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_address <= main_genericstandalone_rtio_core_sed_record43_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_data <= main_genericstandalone_rtio_core_sed_record43_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record63_rec_valid <= main_genericstandalone_rtio_core_sed_record47_rec_valid;
			main_genericstandalone_rtio_core_sed_record63_rec_seqn <= main_genericstandalone_rtio_core_sed_record47_rec_seqn;
			main_genericstandalone_rtio_core_sed_record63_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record47_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record63_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record47_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record47_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record47_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_address <= main_genericstandalone_rtio_core_sed_record47_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_data <= main_genericstandalone_rtio_core_sed_record47_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record59_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference27;
		main_genericstandalone_rtio_core_sed_record63_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record43_rec_valid), main_genericstandalone_rtio_core_sed_record43_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record47_rec_valid), main_genericstandalone_rtio_core_sed_record47_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record59_rec_valid <= main_genericstandalone_rtio_core_sed_record43_rec_valid;
			main_genericstandalone_rtio_core_sed_record59_rec_seqn <= main_genericstandalone_rtio_core_sed_record43_rec_seqn;
			main_genericstandalone_rtio_core_sed_record59_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record43_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record43_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record43_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record43_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_address <= main_genericstandalone_rtio_core_sed_record43_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_data <= main_genericstandalone_rtio_core_sed_record43_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record63_rec_valid <= main_genericstandalone_rtio_core_sed_record47_rec_valid;
			main_genericstandalone_rtio_core_sed_record63_rec_seqn <= main_genericstandalone_rtio_core_sed_record47_rec_seqn;
			main_genericstandalone_rtio_core_sed_record63_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record47_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record63_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record47_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record47_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record47_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_address <= main_genericstandalone_rtio_core_sed_record47_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_data <= main_genericstandalone_rtio_core_sed_record47_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record59_rec_valid <= main_genericstandalone_rtio_core_sed_record47_rec_valid;
			main_genericstandalone_rtio_core_sed_record59_rec_seqn <= main_genericstandalone_rtio_core_sed_record47_rec_seqn;
			main_genericstandalone_rtio_core_sed_record59_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record47_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record47_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record47_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record47_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_address <= main_genericstandalone_rtio_core_sed_record47_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record59_rec_payload_data <= main_genericstandalone_rtio_core_sed_record47_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record63_rec_valid <= main_genericstandalone_rtio_core_sed_record43_rec_valid;
			main_genericstandalone_rtio_core_sed_record63_rec_seqn <= main_genericstandalone_rtio_core_sed_record43_rec_seqn;
			main_genericstandalone_rtio_core_sed_record63_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record43_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record63_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record43_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record43_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record43_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_address <= main_genericstandalone_rtio_core_sed_record43_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record63_rec_payload_data <= main_genericstandalone_rtio_core_sed_record43_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record50_rec_valid), main_genericstandalone_rtio_core_sed_record50_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record52_rec_valid), main_genericstandalone_rtio_core_sed_record52_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record50_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record50_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record52_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record52_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record50_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record52_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record50_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record50_rec_seqn < main_genericstandalone_rtio_core_sed_record52_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record66_rec_valid <= main_genericstandalone_rtio_core_sed_record52_rec_valid;
			main_genericstandalone_rtio_core_sed_record66_rec_seqn <= main_genericstandalone_rtio_core_sed_record52_rec_seqn;
			main_genericstandalone_rtio_core_sed_record66_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record52_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record52_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_address <= main_genericstandalone_rtio_core_sed_record52_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_data <= main_genericstandalone_rtio_core_sed_record52_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record68_rec_valid <= main_genericstandalone_rtio_core_sed_record50_rec_valid;
			main_genericstandalone_rtio_core_sed_record68_rec_seqn <= main_genericstandalone_rtio_core_sed_record50_rec_seqn;
			main_genericstandalone_rtio_core_sed_record68_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record50_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record50_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_address <= main_genericstandalone_rtio_core_sed_record50_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_data <= main_genericstandalone_rtio_core_sed_record50_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record66_rec_valid <= main_genericstandalone_rtio_core_sed_record50_rec_valid;
			main_genericstandalone_rtio_core_sed_record66_rec_seqn <= main_genericstandalone_rtio_core_sed_record50_rec_seqn;
			main_genericstandalone_rtio_core_sed_record66_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record50_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record50_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_address <= main_genericstandalone_rtio_core_sed_record50_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_data <= main_genericstandalone_rtio_core_sed_record50_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record68_rec_valid <= main_genericstandalone_rtio_core_sed_record52_rec_valid;
			main_genericstandalone_rtio_core_sed_record68_rec_seqn <= main_genericstandalone_rtio_core_sed_record52_rec_seqn;
			main_genericstandalone_rtio_core_sed_record68_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record52_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record52_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_address <= main_genericstandalone_rtio_core_sed_record52_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_data <= main_genericstandalone_rtio_core_sed_record52_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record66_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference28;
		main_genericstandalone_rtio_core_sed_record68_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record50_rec_valid), main_genericstandalone_rtio_core_sed_record50_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record52_rec_valid), main_genericstandalone_rtio_core_sed_record52_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record66_rec_valid <= main_genericstandalone_rtio_core_sed_record50_rec_valid;
			main_genericstandalone_rtio_core_sed_record66_rec_seqn <= main_genericstandalone_rtio_core_sed_record50_rec_seqn;
			main_genericstandalone_rtio_core_sed_record66_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record50_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record50_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_address <= main_genericstandalone_rtio_core_sed_record50_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_data <= main_genericstandalone_rtio_core_sed_record50_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record68_rec_valid <= main_genericstandalone_rtio_core_sed_record52_rec_valid;
			main_genericstandalone_rtio_core_sed_record68_rec_seqn <= main_genericstandalone_rtio_core_sed_record52_rec_seqn;
			main_genericstandalone_rtio_core_sed_record68_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record52_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record52_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_address <= main_genericstandalone_rtio_core_sed_record52_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_data <= main_genericstandalone_rtio_core_sed_record52_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record66_rec_valid <= main_genericstandalone_rtio_core_sed_record52_rec_valid;
			main_genericstandalone_rtio_core_sed_record66_rec_seqn <= main_genericstandalone_rtio_core_sed_record52_rec_seqn;
			main_genericstandalone_rtio_core_sed_record66_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record52_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record52_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record52_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record52_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_address <= main_genericstandalone_rtio_core_sed_record52_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record66_rec_payload_data <= main_genericstandalone_rtio_core_sed_record52_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record68_rec_valid <= main_genericstandalone_rtio_core_sed_record50_rec_valid;
			main_genericstandalone_rtio_core_sed_record68_rec_seqn <= main_genericstandalone_rtio_core_sed_record50_rec_seqn;
			main_genericstandalone_rtio_core_sed_record68_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record50_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record50_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record50_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record50_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_address <= main_genericstandalone_rtio_core_sed_record50_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record68_rec_payload_data <= main_genericstandalone_rtio_core_sed_record50_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record51_rec_valid), main_genericstandalone_rtio_core_sed_record51_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record53_rec_valid), main_genericstandalone_rtio_core_sed_record53_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record51_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record51_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record53_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record53_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record51_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record53_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record51_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record51_rec_seqn < main_genericstandalone_rtio_core_sed_record53_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record67_rec_valid <= main_genericstandalone_rtio_core_sed_record53_rec_valid;
			main_genericstandalone_rtio_core_sed_record67_rec_seqn <= main_genericstandalone_rtio_core_sed_record53_rec_seqn;
			main_genericstandalone_rtio_core_sed_record67_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record53_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record53_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_address <= main_genericstandalone_rtio_core_sed_record53_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_data <= main_genericstandalone_rtio_core_sed_record53_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record69_rec_valid <= main_genericstandalone_rtio_core_sed_record51_rec_valid;
			main_genericstandalone_rtio_core_sed_record69_rec_seqn <= main_genericstandalone_rtio_core_sed_record51_rec_seqn;
			main_genericstandalone_rtio_core_sed_record69_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record51_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record51_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_address <= main_genericstandalone_rtio_core_sed_record51_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_data <= main_genericstandalone_rtio_core_sed_record51_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record67_rec_valid <= main_genericstandalone_rtio_core_sed_record51_rec_valid;
			main_genericstandalone_rtio_core_sed_record67_rec_seqn <= main_genericstandalone_rtio_core_sed_record51_rec_seqn;
			main_genericstandalone_rtio_core_sed_record67_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record51_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record51_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_address <= main_genericstandalone_rtio_core_sed_record51_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_data <= main_genericstandalone_rtio_core_sed_record51_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record69_rec_valid <= main_genericstandalone_rtio_core_sed_record53_rec_valid;
			main_genericstandalone_rtio_core_sed_record69_rec_seqn <= main_genericstandalone_rtio_core_sed_record53_rec_seqn;
			main_genericstandalone_rtio_core_sed_record69_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record53_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record53_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_address <= main_genericstandalone_rtio_core_sed_record53_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_data <= main_genericstandalone_rtio_core_sed_record53_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record67_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference29;
		main_genericstandalone_rtio_core_sed_record69_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record51_rec_valid), main_genericstandalone_rtio_core_sed_record51_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record53_rec_valid), main_genericstandalone_rtio_core_sed_record53_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record67_rec_valid <= main_genericstandalone_rtio_core_sed_record51_rec_valid;
			main_genericstandalone_rtio_core_sed_record67_rec_seqn <= main_genericstandalone_rtio_core_sed_record51_rec_seqn;
			main_genericstandalone_rtio_core_sed_record67_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record51_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record51_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_address <= main_genericstandalone_rtio_core_sed_record51_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_data <= main_genericstandalone_rtio_core_sed_record51_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record69_rec_valid <= main_genericstandalone_rtio_core_sed_record53_rec_valid;
			main_genericstandalone_rtio_core_sed_record69_rec_seqn <= main_genericstandalone_rtio_core_sed_record53_rec_seqn;
			main_genericstandalone_rtio_core_sed_record69_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record53_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record53_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_address <= main_genericstandalone_rtio_core_sed_record53_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_data <= main_genericstandalone_rtio_core_sed_record53_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record67_rec_valid <= main_genericstandalone_rtio_core_sed_record53_rec_valid;
			main_genericstandalone_rtio_core_sed_record67_rec_seqn <= main_genericstandalone_rtio_core_sed_record53_rec_seqn;
			main_genericstandalone_rtio_core_sed_record67_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record53_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record53_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record53_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record53_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_address <= main_genericstandalone_rtio_core_sed_record53_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record67_rec_payload_data <= main_genericstandalone_rtio_core_sed_record53_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record69_rec_valid <= main_genericstandalone_rtio_core_sed_record51_rec_valid;
			main_genericstandalone_rtio_core_sed_record69_rec_seqn <= main_genericstandalone_rtio_core_sed_record51_rec_seqn;
			main_genericstandalone_rtio_core_sed_record69_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record51_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record51_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record51_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record51_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_address <= main_genericstandalone_rtio_core_sed_record51_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record69_rec_payload_data <= main_genericstandalone_rtio_core_sed_record51_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record58_rec_valid), main_genericstandalone_rtio_core_sed_record58_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record60_rec_valid), main_genericstandalone_rtio_core_sed_record60_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record58_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record58_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record60_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record60_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record58_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record60_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record58_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record58_rec_seqn < main_genericstandalone_rtio_core_sed_record60_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record74_rec_valid <= main_genericstandalone_rtio_core_sed_record60_rec_valid;
			main_genericstandalone_rtio_core_sed_record74_rec_seqn <= main_genericstandalone_rtio_core_sed_record60_rec_seqn;
			main_genericstandalone_rtio_core_sed_record74_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record60_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record60_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_address <= main_genericstandalone_rtio_core_sed_record60_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_data <= main_genericstandalone_rtio_core_sed_record60_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record76_rec_valid <= main_genericstandalone_rtio_core_sed_record58_rec_valid;
			main_genericstandalone_rtio_core_sed_record76_rec_seqn <= main_genericstandalone_rtio_core_sed_record58_rec_seqn;
			main_genericstandalone_rtio_core_sed_record76_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record58_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record58_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_address <= main_genericstandalone_rtio_core_sed_record58_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_data <= main_genericstandalone_rtio_core_sed_record58_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record74_rec_valid <= main_genericstandalone_rtio_core_sed_record58_rec_valid;
			main_genericstandalone_rtio_core_sed_record74_rec_seqn <= main_genericstandalone_rtio_core_sed_record58_rec_seqn;
			main_genericstandalone_rtio_core_sed_record74_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record58_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record58_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_address <= main_genericstandalone_rtio_core_sed_record58_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_data <= main_genericstandalone_rtio_core_sed_record58_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record76_rec_valid <= main_genericstandalone_rtio_core_sed_record60_rec_valid;
			main_genericstandalone_rtio_core_sed_record76_rec_seqn <= main_genericstandalone_rtio_core_sed_record60_rec_seqn;
			main_genericstandalone_rtio_core_sed_record76_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record60_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record60_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_address <= main_genericstandalone_rtio_core_sed_record60_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_data <= main_genericstandalone_rtio_core_sed_record60_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record74_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference30;
		main_genericstandalone_rtio_core_sed_record76_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record58_rec_valid), main_genericstandalone_rtio_core_sed_record58_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record60_rec_valid), main_genericstandalone_rtio_core_sed_record60_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record74_rec_valid <= main_genericstandalone_rtio_core_sed_record58_rec_valid;
			main_genericstandalone_rtio_core_sed_record74_rec_seqn <= main_genericstandalone_rtio_core_sed_record58_rec_seqn;
			main_genericstandalone_rtio_core_sed_record74_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record58_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record58_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_address <= main_genericstandalone_rtio_core_sed_record58_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_data <= main_genericstandalone_rtio_core_sed_record58_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record76_rec_valid <= main_genericstandalone_rtio_core_sed_record60_rec_valid;
			main_genericstandalone_rtio_core_sed_record76_rec_seqn <= main_genericstandalone_rtio_core_sed_record60_rec_seqn;
			main_genericstandalone_rtio_core_sed_record76_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record60_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record60_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_address <= main_genericstandalone_rtio_core_sed_record60_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_data <= main_genericstandalone_rtio_core_sed_record60_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record74_rec_valid <= main_genericstandalone_rtio_core_sed_record60_rec_valid;
			main_genericstandalone_rtio_core_sed_record74_rec_seqn <= main_genericstandalone_rtio_core_sed_record60_rec_seqn;
			main_genericstandalone_rtio_core_sed_record74_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record60_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record60_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record60_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record60_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_address <= main_genericstandalone_rtio_core_sed_record60_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record74_rec_payload_data <= main_genericstandalone_rtio_core_sed_record60_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record76_rec_valid <= main_genericstandalone_rtio_core_sed_record58_rec_valid;
			main_genericstandalone_rtio_core_sed_record76_rec_seqn <= main_genericstandalone_rtio_core_sed_record58_rec_seqn;
			main_genericstandalone_rtio_core_sed_record76_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record58_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record58_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record58_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record58_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_address <= main_genericstandalone_rtio_core_sed_record58_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record76_rec_payload_data <= main_genericstandalone_rtio_core_sed_record58_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record59_rec_valid), main_genericstandalone_rtio_core_sed_record59_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record61_rec_valid), main_genericstandalone_rtio_core_sed_record61_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record59_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record59_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record61_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record61_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record59_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record61_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record59_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record59_rec_seqn < main_genericstandalone_rtio_core_sed_record61_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record75_rec_valid <= main_genericstandalone_rtio_core_sed_record61_rec_valid;
			main_genericstandalone_rtio_core_sed_record75_rec_seqn <= main_genericstandalone_rtio_core_sed_record61_rec_seqn;
			main_genericstandalone_rtio_core_sed_record75_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record61_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record61_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_address <= main_genericstandalone_rtio_core_sed_record61_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_data <= main_genericstandalone_rtio_core_sed_record61_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record77_rec_valid <= main_genericstandalone_rtio_core_sed_record59_rec_valid;
			main_genericstandalone_rtio_core_sed_record77_rec_seqn <= main_genericstandalone_rtio_core_sed_record59_rec_seqn;
			main_genericstandalone_rtio_core_sed_record77_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record59_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record59_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_address <= main_genericstandalone_rtio_core_sed_record59_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_data <= main_genericstandalone_rtio_core_sed_record59_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record75_rec_valid <= main_genericstandalone_rtio_core_sed_record59_rec_valid;
			main_genericstandalone_rtio_core_sed_record75_rec_seqn <= main_genericstandalone_rtio_core_sed_record59_rec_seqn;
			main_genericstandalone_rtio_core_sed_record75_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record59_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record59_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_address <= main_genericstandalone_rtio_core_sed_record59_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_data <= main_genericstandalone_rtio_core_sed_record59_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record77_rec_valid <= main_genericstandalone_rtio_core_sed_record61_rec_valid;
			main_genericstandalone_rtio_core_sed_record77_rec_seqn <= main_genericstandalone_rtio_core_sed_record61_rec_seqn;
			main_genericstandalone_rtio_core_sed_record77_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record61_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record61_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_address <= main_genericstandalone_rtio_core_sed_record61_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_data <= main_genericstandalone_rtio_core_sed_record61_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record75_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference31;
		main_genericstandalone_rtio_core_sed_record77_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record59_rec_valid), main_genericstandalone_rtio_core_sed_record59_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record61_rec_valid), main_genericstandalone_rtio_core_sed_record61_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record75_rec_valid <= main_genericstandalone_rtio_core_sed_record59_rec_valid;
			main_genericstandalone_rtio_core_sed_record75_rec_seqn <= main_genericstandalone_rtio_core_sed_record59_rec_seqn;
			main_genericstandalone_rtio_core_sed_record75_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record59_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record59_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_address <= main_genericstandalone_rtio_core_sed_record59_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_data <= main_genericstandalone_rtio_core_sed_record59_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record77_rec_valid <= main_genericstandalone_rtio_core_sed_record61_rec_valid;
			main_genericstandalone_rtio_core_sed_record77_rec_seqn <= main_genericstandalone_rtio_core_sed_record61_rec_seqn;
			main_genericstandalone_rtio_core_sed_record77_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record61_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record61_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_address <= main_genericstandalone_rtio_core_sed_record61_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_data <= main_genericstandalone_rtio_core_sed_record61_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record75_rec_valid <= main_genericstandalone_rtio_core_sed_record61_rec_valid;
			main_genericstandalone_rtio_core_sed_record75_rec_seqn <= main_genericstandalone_rtio_core_sed_record61_rec_seqn;
			main_genericstandalone_rtio_core_sed_record75_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record61_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record61_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record61_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record61_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_address <= main_genericstandalone_rtio_core_sed_record61_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record75_rec_payload_data <= main_genericstandalone_rtio_core_sed_record61_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record77_rec_valid <= main_genericstandalone_rtio_core_sed_record59_rec_valid;
			main_genericstandalone_rtio_core_sed_record77_rec_seqn <= main_genericstandalone_rtio_core_sed_record59_rec_seqn;
			main_genericstandalone_rtio_core_sed_record77_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record59_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record59_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record59_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record59_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_address <= main_genericstandalone_rtio_core_sed_record59_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record77_rec_payload_data <= main_genericstandalone_rtio_core_sed_record59_rec_payload_data;
		end
	end
	main_genericstandalone_rtio_core_sed_record64_rec_valid <= main_genericstandalone_rtio_core_sed_record48_rec_valid;
	main_genericstandalone_rtio_core_sed_record64_rec_seqn <= main_genericstandalone_rtio_core_sed_record48_rec_seqn;
	main_genericstandalone_rtio_core_sed_record64_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record48_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record64_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record48_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record64_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record48_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record64_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record48_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record64_rec_payload_address <= main_genericstandalone_rtio_core_sed_record48_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record64_rec_payload_data <= main_genericstandalone_rtio_core_sed_record48_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record65_rec_valid <= main_genericstandalone_rtio_core_sed_record49_rec_valid;
	main_genericstandalone_rtio_core_sed_record65_rec_seqn <= main_genericstandalone_rtio_core_sed_record49_rec_seqn;
	main_genericstandalone_rtio_core_sed_record65_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record49_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record65_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record49_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record65_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record49_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record65_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record49_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record65_rec_payload_address <= main_genericstandalone_rtio_core_sed_record49_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record65_rec_payload_data <= main_genericstandalone_rtio_core_sed_record49_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record70_rec_valid <= main_genericstandalone_rtio_core_sed_record54_rec_valid;
	main_genericstandalone_rtio_core_sed_record70_rec_seqn <= main_genericstandalone_rtio_core_sed_record54_rec_seqn;
	main_genericstandalone_rtio_core_sed_record70_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record54_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record70_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record54_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record70_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record54_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record70_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record54_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record70_rec_payload_address <= main_genericstandalone_rtio_core_sed_record54_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record70_rec_payload_data <= main_genericstandalone_rtio_core_sed_record54_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record71_rec_valid <= main_genericstandalone_rtio_core_sed_record55_rec_valid;
	main_genericstandalone_rtio_core_sed_record71_rec_seqn <= main_genericstandalone_rtio_core_sed_record55_rec_seqn;
	main_genericstandalone_rtio_core_sed_record71_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record55_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record71_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record55_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record71_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record55_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record71_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record55_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record71_rec_payload_address <= main_genericstandalone_rtio_core_sed_record55_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record71_rec_payload_data <= main_genericstandalone_rtio_core_sed_record55_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record72_rec_valid <= main_genericstandalone_rtio_core_sed_record56_rec_valid;
	main_genericstandalone_rtio_core_sed_record72_rec_seqn <= main_genericstandalone_rtio_core_sed_record56_rec_seqn;
	main_genericstandalone_rtio_core_sed_record72_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record56_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record72_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record56_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record72_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record56_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record72_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record56_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record72_rec_payload_address <= main_genericstandalone_rtio_core_sed_record56_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record72_rec_payload_data <= main_genericstandalone_rtio_core_sed_record56_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record73_rec_valid <= main_genericstandalone_rtio_core_sed_record57_rec_valid;
	main_genericstandalone_rtio_core_sed_record73_rec_seqn <= main_genericstandalone_rtio_core_sed_record57_rec_seqn;
	main_genericstandalone_rtio_core_sed_record73_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record57_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record73_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record57_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record73_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record57_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record73_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record57_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record73_rec_payload_address <= main_genericstandalone_rtio_core_sed_record57_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record73_rec_payload_data <= main_genericstandalone_rtio_core_sed_record57_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record78_rec_valid <= main_genericstandalone_rtio_core_sed_record62_rec_valid;
	main_genericstandalone_rtio_core_sed_record78_rec_seqn <= main_genericstandalone_rtio_core_sed_record62_rec_seqn;
	main_genericstandalone_rtio_core_sed_record78_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record62_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record78_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record62_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record78_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record62_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record78_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record62_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record78_rec_payload_address <= main_genericstandalone_rtio_core_sed_record62_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record78_rec_payload_data <= main_genericstandalone_rtio_core_sed_record62_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record79_rec_valid <= main_genericstandalone_rtio_core_sed_record63_rec_valid;
	main_genericstandalone_rtio_core_sed_record79_rec_seqn <= main_genericstandalone_rtio_core_sed_record63_rec_seqn;
	main_genericstandalone_rtio_core_sed_record79_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record63_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record79_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record63_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record79_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record63_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record79_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record63_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record79_rec_payload_address <= main_genericstandalone_rtio_core_sed_record63_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record79_rec_payload_data <= main_genericstandalone_rtio_core_sed_record63_rec_payload_data;
	if (({(~main_genericstandalone_rtio_core_sed_record65_rec_valid), main_genericstandalone_rtio_core_sed_record65_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record66_rec_valid), main_genericstandalone_rtio_core_sed_record66_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record65_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record65_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record66_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record66_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record65_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record66_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record65_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record65_rec_seqn < main_genericstandalone_rtio_core_sed_record66_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record81_rec_valid <= main_genericstandalone_rtio_core_sed_record66_rec_valid;
			main_genericstandalone_rtio_core_sed_record81_rec_seqn <= main_genericstandalone_rtio_core_sed_record66_rec_seqn;
			main_genericstandalone_rtio_core_sed_record81_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record66_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record66_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_address <= main_genericstandalone_rtio_core_sed_record66_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_data <= main_genericstandalone_rtio_core_sed_record66_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record82_rec_valid <= main_genericstandalone_rtio_core_sed_record65_rec_valid;
			main_genericstandalone_rtio_core_sed_record82_rec_seqn <= main_genericstandalone_rtio_core_sed_record65_rec_seqn;
			main_genericstandalone_rtio_core_sed_record82_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record65_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record65_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record65_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record65_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_address <= main_genericstandalone_rtio_core_sed_record65_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_data <= main_genericstandalone_rtio_core_sed_record65_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record81_rec_valid <= main_genericstandalone_rtio_core_sed_record65_rec_valid;
			main_genericstandalone_rtio_core_sed_record81_rec_seqn <= main_genericstandalone_rtio_core_sed_record65_rec_seqn;
			main_genericstandalone_rtio_core_sed_record81_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record65_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record65_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record65_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record65_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_address <= main_genericstandalone_rtio_core_sed_record65_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_data <= main_genericstandalone_rtio_core_sed_record65_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record82_rec_valid <= main_genericstandalone_rtio_core_sed_record66_rec_valid;
			main_genericstandalone_rtio_core_sed_record82_rec_seqn <= main_genericstandalone_rtio_core_sed_record66_rec_seqn;
			main_genericstandalone_rtio_core_sed_record82_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record66_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record66_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_address <= main_genericstandalone_rtio_core_sed_record66_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_data <= main_genericstandalone_rtio_core_sed_record66_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record81_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference32;
		main_genericstandalone_rtio_core_sed_record82_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record65_rec_valid), main_genericstandalone_rtio_core_sed_record65_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record66_rec_valid), main_genericstandalone_rtio_core_sed_record66_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record81_rec_valid <= main_genericstandalone_rtio_core_sed_record65_rec_valid;
			main_genericstandalone_rtio_core_sed_record81_rec_seqn <= main_genericstandalone_rtio_core_sed_record65_rec_seqn;
			main_genericstandalone_rtio_core_sed_record81_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record65_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record65_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record65_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record65_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_address <= main_genericstandalone_rtio_core_sed_record65_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_data <= main_genericstandalone_rtio_core_sed_record65_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record82_rec_valid <= main_genericstandalone_rtio_core_sed_record66_rec_valid;
			main_genericstandalone_rtio_core_sed_record82_rec_seqn <= main_genericstandalone_rtio_core_sed_record66_rec_seqn;
			main_genericstandalone_rtio_core_sed_record82_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record66_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record66_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_address <= main_genericstandalone_rtio_core_sed_record66_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_data <= main_genericstandalone_rtio_core_sed_record66_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record81_rec_valid <= main_genericstandalone_rtio_core_sed_record66_rec_valid;
			main_genericstandalone_rtio_core_sed_record81_rec_seqn <= main_genericstandalone_rtio_core_sed_record66_rec_seqn;
			main_genericstandalone_rtio_core_sed_record81_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record66_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record66_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record66_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record66_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_address <= main_genericstandalone_rtio_core_sed_record66_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record81_rec_payload_data <= main_genericstandalone_rtio_core_sed_record66_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record82_rec_valid <= main_genericstandalone_rtio_core_sed_record65_rec_valid;
			main_genericstandalone_rtio_core_sed_record82_rec_seqn <= main_genericstandalone_rtio_core_sed_record65_rec_seqn;
			main_genericstandalone_rtio_core_sed_record82_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record65_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record65_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record65_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record65_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_address <= main_genericstandalone_rtio_core_sed_record65_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record82_rec_payload_data <= main_genericstandalone_rtio_core_sed_record65_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record67_rec_valid), main_genericstandalone_rtio_core_sed_record67_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record68_rec_valid), main_genericstandalone_rtio_core_sed_record68_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record67_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record67_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record68_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record68_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record67_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record68_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record67_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record67_rec_seqn < main_genericstandalone_rtio_core_sed_record68_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record83_rec_valid <= main_genericstandalone_rtio_core_sed_record68_rec_valid;
			main_genericstandalone_rtio_core_sed_record83_rec_seqn <= main_genericstandalone_rtio_core_sed_record68_rec_seqn;
			main_genericstandalone_rtio_core_sed_record83_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record68_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record68_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_address <= main_genericstandalone_rtio_core_sed_record68_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_data <= main_genericstandalone_rtio_core_sed_record68_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record84_rec_valid <= main_genericstandalone_rtio_core_sed_record67_rec_valid;
			main_genericstandalone_rtio_core_sed_record84_rec_seqn <= main_genericstandalone_rtio_core_sed_record67_rec_seqn;
			main_genericstandalone_rtio_core_sed_record84_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record67_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record67_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_address <= main_genericstandalone_rtio_core_sed_record67_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_data <= main_genericstandalone_rtio_core_sed_record67_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record83_rec_valid <= main_genericstandalone_rtio_core_sed_record67_rec_valid;
			main_genericstandalone_rtio_core_sed_record83_rec_seqn <= main_genericstandalone_rtio_core_sed_record67_rec_seqn;
			main_genericstandalone_rtio_core_sed_record83_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record67_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record67_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_address <= main_genericstandalone_rtio_core_sed_record67_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_data <= main_genericstandalone_rtio_core_sed_record67_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record84_rec_valid <= main_genericstandalone_rtio_core_sed_record68_rec_valid;
			main_genericstandalone_rtio_core_sed_record84_rec_seqn <= main_genericstandalone_rtio_core_sed_record68_rec_seqn;
			main_genericstandalone_rtio_core_sed_record84_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record68_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record68_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_address <= main_genericstandalone_rtio_core_sed_record68_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_data <= main_genericstandalone_rtio_core_sed_record68_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record83_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference33;
		main_genericstandalone_rtio_core_sed_record84_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record67_rec_valid), main_genericstandalone_rtio_core_sed_record67_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record68_rec_valid), main_genericstandalone_rtio_core_sed_record68_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record83_rec_valid <= main_genericstandalone_rtio_core_sed_record67_rec_valid;
			main_genericstandalone_rtio_core_sed_record83_rec_seqn <= main_genericstandalone_rtio_core_sed_record67_rec_seqn;
			main_genericstandalone_rtio_core_sed_record83_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record67_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record67_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_address <= main_genericstandalone_rtio_core_sed_record67_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_data <= main_genericstandalone_rtio_core_sed_record67_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record84_rec_valid <= main_genericstandalone_rtio_core_sed_record68_rec_valid;
			main_genericstandalone_rtio_core_sed_record84_rec_seqn <= main_genericstandalone_rtio_core_sed_record68_rec_seqn;
			main_genericstandalone_rtio_core_sed_record84_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record68_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record68_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_address <= main_genericstandalone_rtio_core_sed_record68_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_data <= main_genericstandalone_rtio_core_sed_record68_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record83_rec_valid <= main_genericstandalone_rtio_core_sed_record68_rec_valid;
			main_genericstandalone_rtio_core_sed_record83_rec_seqn <= main_genericstandalone_rtio_core_sed_record68_rec_seqn;
			main_genericstandalone_rtio_core_sed_record83_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record68_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record68_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record68_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record68_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_address <= main_genericstandalone_rtio_core_sed_record68_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record83_rec_payload_data <= main_genericstandalone_rtio_core_sed_record68_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record84_rec_valid <= main_genericstandalone_rtio_core_sed_record67_rec_valid;
			main_genericstandalone_rtio_core_sed_record84_rec_seqn <= main_genericstandalone_rtio_core_sed_record67_rec_seqn;
			main_genericstandalone_rtio_core_sed_record84_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record67_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record67_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record67_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record67_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_address <= main_genericstandalone_rtio_core_sed_record67_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record84_rec_payload_data <= main_genericstandalone_rtio_core_sed_record67_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record69_rec_valid), main_genericstandalone_rtio_core_sed_record69_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record70_rec_valid), main_genericstandalone_rtio_core_sed_record70_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record69_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record69_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record70_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record70_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record69_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record70_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record69_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record69_rec_seqn < main_genericstandalone_rtio_core_sed_record70_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record85_rec_valid <= main_genericstandalone_rtio_core_sed_record70_rec_valid;
			main_genericstandalone_rtio_core_sed_record85_rec_seqn <= main_genericstandalone_rtio_core_sed_record70_rec_seqn;
			main_genericstandalone_rtio_core_sed_record85_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record70_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record70_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record70_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record70_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_address <= main_genericstandalone_rtio_core_sed_record70_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_data <= main_genericstandalone_rtio_core_sed_record70_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record86_rec_valid <= main_genericstandalone_rtio_core_sed_record69_rec_valid;
			main_genericstandalone_rtio_core_sed_record86_rec_seqn <= main_genericstandalone_rtio_core_sed_record69_rec_seqn;
			main_genericstandalone_rtio_core_sed_record86_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record69_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record69_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_address <= main_genericstandalone_rtio_core_sed_record69_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_data <= main_genericstandalone_rtio_core_sed_record69_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record85_rec_valid <= main_genericstandalone_rtio_core_sed_record69_rec_valid;
			main_genericstandalone_rtio_core_sed_record85_rec_seqn <= main_genericstandalone_rtio_core_sed_record69_rec_seqn;
			main_genericstandalone_rtio_core_sed_record85_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record69_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record69_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_address <= main_genericstandalone_rtio_core_sed_record69_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_data <= main_genericstandalone_rtio_core_sed_record69_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record86_rec_valid <= main_genericstandalone_rtio_core_sed_record70_rec_valid;
			main_genericstandalone_rtio_core_sed_record86_rec_seqn <= main_genericstandalone_rtio_core_sed_record70_rec_seqn;
			main_genericstandalone_rtio_core_sed_record86_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record70_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record70_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record70_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record70_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_address <= main_genericstandalone_rtio_core_sed_record70_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_data <= main_genericstandalone_rtio_core_sed_record70_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record85_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference34;
		main_genericstandalone_rtio_core_sed_record86_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record69_rec_valid), main_genericstandalone_rtio_core_sed_record69_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record70_rec_valid), main_genericstandalone_rtio_core_sed_record70_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record85_rec_valid <= main_genericstandalone_rtio_core_sed_record69_rec_valid;
			main_genericstandalone_rtio_core_sed_record85_rec_seqn <= main_genericstandalone_rtio_core_sed_record69_rec_seqn;
			main_genericstandalone_rtio_core_sed_record85_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record69_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record69_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_address <= main_genericstandalone_rtio_core_sed_record69_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_data <= main_genericstandalone_rtio_core_sed_record69_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record86_rec_valid <= main_genericstandalone_rtio_core_sed_record70_rec_valid;
			main_genericstandalone_rtio_core_sed_record86_rec_seqn <= main_genericstandalone_rtio_core_sed_record70_rec_seqn;
			main_genericstandalone_rtio_core_sed_record86_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record70_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record70_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record70_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record70_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_address <= main_genericstandalone_rtio_core_sed_record70_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_data <= main_genericstandalone_rtio_core_sed_record70_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record85_rec_valid <= main_genericstandalone_rtio_core_sed_record70_rec_valid;
			main_genericstandalone_rtio_core_sed_record85_rec_seqn <= main_genericstandalone_rtio_core_sed_record70_rec_seqn;
			main_genericstandalone_rtio_core_sed_record85_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record70_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record70_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record70_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record70_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_address <= main_genericstandalone_rtio_core_sed_record70_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record85_rec_payload_data <= main_genericstandalone_rtio_core_sed_record70_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record86_rec_valid <= main_genericstandalone_rtio_core_sed_record69_rec_valid;
			main_genericstandalone_rtio_core_sed_record86_rec_seqn <= main_genericstandalone_rtio_core_sed_record69_rec_seqn;
			main_genericstandalone_rtio_core_sed_record86_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record69_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record69_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record69_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record69_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_address <= main_genericstandalone_rtio_core_sed_record69_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record86_rec_payload_data <= main_genericstandalone_rtio_core_sed_record69_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record73_rec_valid), main_genericstandalone_rtio_core_sed_record73_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record74_rec_valid), main_genericstandalone_rtio_core_sed_record74_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record73_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record73_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record74_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record74_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record73_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record74_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record73_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record73_rec_seqn < main_genericstandalone_rtio_core_sed_record74_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record89_rec_valid <= main_genericstandalone_rtio_core_sed_record74_rec_valid;
			main_genericstandalone_rtio_core_sed_record89_rec_seqn <= main_genericstandalone_rtio_core_sed_record74_rec_seqn;
			main_genericstandalone_rtio_core_sed_record89_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record74_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record74_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_address <= main_genericstandalone_rtio_core_sed_record74_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_data <= main_genericstandalone_rtio_core_sed_record74_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record90_rec_valid <= main_genericstandalone_rtio_core_sed_record73_rec_valid;
			main_genericstandalone_rtio_core_sed_record90_rec_seqn <= main_genericstandalone_rtio_core_sed_record73_rec_seqn;
			main_genericstandalone_rtio_core_sed_record90_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record73_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record73_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record73_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record73_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_address <= main_genericstandalone_rtio_core_sed_record73_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_data <= main_genericstandalone_rtio_core_sed_record73_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record89_rec_valid <= main_genericstandalone_rtio_core_sed_record73_rec_valid;
			main_genericstandalone_rtio_core_sed_record89_rec_seqn <= main_genericstandalone_rtio_core_sed_record73_rec_seqn;
			main_genericstandalone_rtio_core_sed_record89_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record73_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record73_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record73_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record73_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_address <= main_genericstandalone_rtio_core_sed_record73_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_data <= main_genericstandalone_rtio_core_sed_record73_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record90_rec_valid <= main_genericstandalone_rtio_core_sed_record74_rec_valid;
			main_genericstandalone_rtio_core_sed_record90_rec_seqn <= main_genericstandalone_rtio_core_sed_record74_rec_seqn;
			main_genericstandalone_rtio_core_sed_record90_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record74_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record74_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_address <= main_genericstandalone_rtio_core_sed_record74_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_data <= main_genericstandalone_rtio_core_sed_record74_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record89_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference35;
		main_genericstandalone_rtio_core_sed_record90_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record73_rec_valid), main_genericstandalone_rtio_core_sed_record73_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record74_rec_valid), main_genericstandalone_rtio_core_sed_record74_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record89_rec_valid <= main_genericstandalone_rtio_core_sed_record73_rec_valid;
			main_genericstandalone_rtio_core_sed_record89_rec_seqn <= main_genericstandalone_rtio_core_sed_record73_rec_seqn;
			main_genericstandalone_rtio_core_sed_record89_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record73_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record73_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record73_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record73_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_address <= main_genericstandalone_rtio_core_sed_record73_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_data <= main_genericstandalone_rtio_core_sed_record73_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record90_rec_valid <= main_genericstandalone_rtio_core_sed_record74_rec_valid;
			main_genericstandalone_rtio_core_sed_record90_rec_seqn <= main_genericstandalone_rtio_core_sed_record74_rec_seqn;
			main_genericstandalone_rtio_core_sed_record90_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record74_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record74_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_address <= main_genericstandalone_rtio_core_sed_record74_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_data <= main_genericstandalone_rtio_core_sed_record74_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record89_rec_valid <= main_genericstandalone_rtio_core_sed_record74_rec_valid;
			main_genericstandalone_rtio_core_sed_record89_rec_seqn <= main_genericstandalone_rtio_core_sed_record74_rec_seqn;
			main_genericstandalone_rtio_core_sed_record89_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record74_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record74_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record74_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record74_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_address <= main_genericstandalone_rtio_core_sed_record74_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record89_rec_payload_data <= main_genericstandalone_rtio_core_sed_record74_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record90_rec_valid <= main_genericstandalone_rtio_core_sed_record73_rec_valid;
			main_genericstandalone_rtio_core_sed_record90_rec_seqn <= main_genericstandalone_rtio_core_sed_record73_rec_seqn;
			main_genericstandalone_rtio_core_sed_record90_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record73_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record73_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record73_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record73_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_address <= main_genericstandalone_rtio_core_sed_record73_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record90_rec_payload_data <= main_genericstandalone_rtio_core_sed_record73_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record75_rec_valid), main_genericstandalone_rtio_core_sed_record75_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record76_rec_valid), main_genericstandalone_rtio_core_sed_record76_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record75_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record75_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record76_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record76_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record75_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record76_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record75_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record75_rec_seqn < main_genericstandalone_rtio_core_sed_record76_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record91_rec_valid <= main_genericstandalone_rtio_core_sed_record76_rec_valid;
			main_genericstandalone_rtio_core_sed_record91_rec_seqn <= main_genericstandalone_rtio_core_sed_record76_rec_seqn;
			main_genericstandalone_rtio_core_sed_record91_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record76_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record76_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_address <= main_genericstandalone_rtio_core_sed_record76_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_data <= main_genericstandalone_rtio_core_sed_record76_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record92_rec_valid <= main_genericstandalone_rtio_core_sed_record75_rec_valid;
			main_genericstandalone_rtio_core_sed_record92_rec_seqn <= main_genericstandalone_rtio_core_sed_record75_rec_seqn;
			main_genericstandalone_rtio_core_sed_record92_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record75_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record75_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_address <= main_genericstandalone_rtio_core_sed_record75_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_data <= main_genericstandalone_rtio_core_sed_record75_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record91_rec_valid <= main_genericstandalone_rtio_core_sed_record75_rec_valid;
			main_genericstandalone_rtio_core_sed_record91_rec_seqn <= main_genericstandalone_rtio_core_sed_record75_rec_seqn;
			main_genericstandalone_rtio_core_sed_record91_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record75_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record75_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_address <= main_genericstandalone_rtio_core_sed_record75_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_data <= main_genericstandalone_rtio_core_sed_record75_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record92_rec_valid <= main_genericstandalone_rtio_core_sed_record76_rec_valid;
			main_genericstandalone_rtio_core_sed_record92_rec_seqn <= main_genericstandalone_rtio_core_sed_record76_rec_seqn;
			main_genericstandalone_rtio_core_sed_record92_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record76_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record76_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_address <= main_genericstandalone_rtio_core_sed_record76_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_data <= main_genericstandalone_rtio_core_sed_record76_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record91_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference36;
		main_genericstandalone_rtio_core_sed_record92_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record75_rec_valid), main_genericstandalone_rtio_core_sed_record75_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record76_rec_valid), main_genericstandalone_rtio_core_sed_record76_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record91_rec_valid <= main_genericstandalone_rtio_core_sed_record75_rec_valid;
			main_genericstandalone_rtio_core_sed_record91_rec_seqn <= main_genericstandalone_rtio_core_sed_record75_rec_seqn;
			main_genericstandalone_rtio_core_sed_record91_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record75_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record75_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_address <= main_genericstandalone_rtio_core_sed_record75_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_data <= main_genericstandalone_rtio_core_sed_record75_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record92_rec_valid <= main_genericstandalone_rtio_core_sed_record76_rec_valid;
			main_genericstandalone_rtio_core_sed_record92_rec_seqn <= main_genericstandalone_rtio_core_sed_record76_rec_seqn;
			main_genericstandalone_rtio_core_sed_record92_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record76_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record76_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_address <= main_genericstandalone_rtio_core_sed_record76_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_data <= main_genericstandalone_rtio_core_sed_record76_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record91_rec_valid <= main_genericstandalone_rtio_core_sed_record76_rec_valid;
			main_genericstandalone_rtio_core_sed_record91_rec_seqn <= main_genericstandalone_rtio_core_sed_record76_rec_seqn;
			main_genericstandalone_rtio_core_sed_record91_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record76_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record76_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record76_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record76_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_address <= main_genericstandalone_rtio_core_sed_record76_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record91_rec_payload_data <= main_genericstandalone_rtio_core_sed_record76_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record92_rec_valid <= main_genericstandalone_rtio_core_sed_record75_rec_valid;
			main_genericstandalone_rtio_core_sed_record92_rec_seqn <= main_genericstandalone_rtio_core_sed_record75_rec_seqn;
			main_genericstandalone_rtio_core_sed_record92_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record75_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record75_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record75_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record75_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_address <= main_genericstandalone_rtio_core_sed_record75_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record92_rec_payload_data <= main_genericstandalone_rtio_core_sed_record75_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record77_rec_valid), main_genericstandalone_rtio_core_sed_record77_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record78_rec_valid), main_genericstandalone_rtio_core_sed_record78_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record77_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record77_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record78_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record78_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record77_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record78_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record77_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record77_rec_seqn < main_genericstandalone_rtio_core_sed_record78_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record93_rec_valid <= main_genericstandalone_rtio_core_sed_record78_rec_valid;
			main_genericstandalone_rtio_core_sed_record93_rec_seqn <= main_genericstandalone_rtio_core_sed_record78_rec_seqn;
			main_genericstandalone_rtio_core_sed_record93_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record78_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record78_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record78_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record78_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_address <= main_genericstandalone_rtio_core_sed_record78_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_data <= main_genericstandalone_rtio_core_sed_record78_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record94_rec_valid <= main_genericstandalone_rtio_core_sed_record77_rec_valid;
			main_genericstandalone_rtio_core_sed_record94_rec_seqn <= main_genericstandalone_rtio_core_sed_record77_rec_seqn;
			main_genericstandalone_rtio_core_sed_record94_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record77_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record77_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_address <= main_genericstandalone_rtio_core_sed_record77_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_data <= main_genericstandalone_rtio_core_sed_record77_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record93_rec_valid <= main_genericstandalone_rtio_core_sed_record77_rec_valid;
			main_genericstandalone_rtio_core_sed_record93_rec_seqn <= main_genericstandalone_rtio_core_sed_record77_rec_seqn;
			main_genericstandalone_rtio_core_sed_record93_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record77_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record77_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_address <= main_genericstandalone_rtio_core_sed_record77_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_data <= main_genericstandalone_rtio_core_sed_record77_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record94_rec_valid <= main_genericstandalone_rtio_core_sed_record78_rec_valid;
			main_genericstandalone_rtio_core_sed_record94_rec_seqn <= main_genericstandalone_rtio_core_sed_record78_rec_seqn;
			main_genericstandalone_rtio_core_sed_record94_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record78_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record78_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record78_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record78_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_address <= main_genericstandalone_rtio_core_sed_record78_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_data <= main_genericstandalone_rtio_core_sed_record78_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record93_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference37;
		main_genericstandalone_rtio_core_sed_record94_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record77_rec_valid), main_genericstandalone_rtio_core_sed_record77_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record78_rec_valid), main_genericstandalone_rtio_core_sed_record78_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record93_rec_valid <= main_genericstandalone_rtio_core_sed_record77_rec_valid;
			main_genericstandalone_rtio_core_sed_record93_rec_seqn <= main_genericstandalone_rtio_core_sed_record77_rec_seqn;
			main_genericstandalone_rtio_core_sed_record93_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record77_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record77_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_address <= main_genericstandalone_rtio_core_sed_record77_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_data <= main_genericstandalone_rtio_core_sed_record77_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record94_rec_valid <= main_genericstandalone_rtio_core_sed_record78_rec_valid;
			main_genericstandalone_rtio_core_sed_record94_rec_seqn <= main_genericstandalone_rtio_core_sed_record78_rec_seqn;
			main_genericstandalone_rtio_core_sed_record94_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record78_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record78_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record78_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record78_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_address <= main_genericstandalone_rtio_core_sed_record78_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_data <= main_genericstandalone_rtio_core_sed_record78_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record93_rec_valid <= main_genericstandalone_rtio_core_sed_record78_rec_valid;
			main_genericstandalone_rtio_core_sed_record93_rec_seqn <= main_genericstandalone_rtio_core_sed_record78_rec_seqn;
			main_genericstandalone_rtio_core_sed_record93_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record78_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record78_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record78_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record78_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_address <= main_genericstandalone_rtio_core_sed_record78_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record93_rec_payload_data <= main_genericstandalone_rtio_core_sed_record78_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record94_rec_valid <= main_genericstandalone_rtio_core_sed_record77_rec_valid;
			main_genericstandalone_rtio_core_sed_record94_rec_seqn <= main_genericstandalone_rtio_core_sed_record77_rec_seqn;
			main_genericstandalone_rtio_core_sed_record94_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record77_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record77_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record77_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record77_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_address <= main_genericstandalone_rtio_core_sed_record77_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record94_rec_payload_data <= main_genericstandalone_rtio_core_sed_record77_rec_payload_data;
		end
	end
	main_genericstandalone_rtio_core_sed_record80_rec_valid <= main_genericstandalone_rtio_core_sed_record64_rec_valid;
	main_genericstandalone_rtio_core_sed_record80_rec_seqn <= main_genericstandalone_rtio_core_sed_record64_rec_seqn;
	main_genericstandalone_rtio_core_sed_record80_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record64_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record80_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record64_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record80_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record64_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record80_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record64_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record80_rec_payload_address <= main_genericstandalone_rtio_core_sed_record64_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record80_rec_payload_data <= main_genericstandalone_rtio_core_sed_record64_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record87_rec_valid <= main_genericstandalone_rtio_core_sed_record71_rec_valid;
	main_genericstandalone_rtio_core_sed_record87_rec_seqn <= main_genericstandalone_rtio_core_sed_record71_rec_seqn;
	main_genericstandalone_rtio_core_sed_record87_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record71_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record87_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record71_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record87_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record71_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record87_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record71_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record87_rec_payload_address <= main_genericstandalone_rtio_core_sed_record71_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record87_rec_payload_data <= main_genericstandalone_rtio_core_sed_record71_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record88_rec_valid <= main_genericstandalone_rtio_core_sed_record72_rec_valid;
	main_genericstandalone_rtio_core_sed_record88_rec_seqn <= main_genericstandalone_rtio_core_sed_record72_rec_seqn;
	main_genericstandalone_rtio_core_sed_record88_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record72_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record88_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record72_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record88_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record72_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record88_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record72_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record88_rec_payload_address <= main_genericstandalone_rtio_core_sed_record72_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record88_rec_payload_data <= main_genericstandalone_rtio_core_sed_record72_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record95_rec_valid <= main_genericstandalone_rtio_core_sed_record79_rec_valid;
	main_genericstandalone_rtio_core_sed_record95_rec_seqn <= main_genericstandalone_rtio_core_sed_record79_rec_seqn;
	main_genericstandalone_rtio_core_sed_record95_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record79_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record95_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record79_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record95_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record79_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record95_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record79_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record95_rec_payload_address <= main_genericstandalone_rtio_core_sed_record79_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record95_rec_payload_data <= main_genericstandalone_rtio_core_sed_record79_rec_payload_data;
	if (({(~main_genericstandalone_rtio_core_sed_record80_rec_valid), main_genericstandalone_rtio_core_sed_record80_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record88_rec_valid), main_genericstandalone_rtio_core_sed_record88_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record80_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record80_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record88_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record88_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record80_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record88_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record80_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record80_rec_seqn < main_genericstandalone_rtio_core_sed_record88_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record96_rec_valid <= main_genericstandalone_rtio_core_sed_record88_rec_valid;
			main_genericstandalone_rtio_core_sed_record96_rec_seqn <= main_genericstandalone_rtio_core_sed_record88_rec_seqn;
			main_genericstandalone_rtio_core_sed_record96_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record88_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record96_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record88_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record88_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record88_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_address <= main_genericstandalone_rtio_core_sed_record88_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_data <= main_genericstandalone_rtio_core_sed_record88_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record104_rec_valid <= main_genericstandalone_rtio_core_sed_record80_rec_valid;
			main_genericstandalone_rtio_core_sed_record104_rec_seqn <= main_genericstandalone_rtio_core_sed_record80_rec_seqn;
			main_genericstandalone_rtio_core_sed_record104_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record80_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record80_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record80_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record80_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_address <= main_genericstandalone_rtio_core_sed_record80_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_data <= main_genericstandalone_rtio_core_sed_record80_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record96_rec_valid <= main_genericstandalone_rtio_core_sed_record80_rec_valid;
			main_genericstandalone_rtio_core_sed_record96_rec_seqn <= main_genericstandalone_rtio_core_sed_record80_rec_seqn;
			main_genericstandalone_rtio_core_sed_record96_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record80_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record96_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record80_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record80_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record80_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_address <= main_genericstandalone_rtio_core_sed_record80_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_data <= main_genericstandalone_rtio_core_sed_record80_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record104_rec_valid <= main_genericstandalone_rtio_core_sed_record88_rec_valid;
			main_genericstandalone_rtio_core_sed_record104_rec_seqn <= main_genericstandalone_rtio_core_sed_record88_rec_seqn;
			main_genericstandalone_rtio_core_sed_record104_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record88_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record88_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record88_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record88_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_address <= main_genericstandalone_rtio_core_sed_record88_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_data <= main_genericstandalone_rtio_core_sed_record88_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record96_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record96_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference38;
		main_genericstandalone_rtio_core_sed_record104_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record80_rec_valid), main_genericstandalone_rtio_core_sed_record80_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record88_rec_valid), main_genericstandalone_rtio_core_sed_record88_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record96_rec_valid <= main_genericstandalone_rtio_core_sed_record80_rec_valid;
			main_genericstandalone_rtio_core_sed_record96_rec_seqn <= main_genericstandalone_rtio_core_sed_record80_rec_seqn;
			main_genericstandalone_rtio_core_sed_record96_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record80_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record96_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record80_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record80_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record80_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_address <= main_genericstandalone_rtio_core_sed_record80_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_data <= main_genericstandalone_rtio_core_sed_record80_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record104_rec_valid <= main_genericstandalone_rtio_core_sed_record88_rec_valid;
			main_genericstandalone_rtio_core_sed_record104_rec_seqn <= main_genericstandalone_rtio_core_sed_record88_rec_seqn;
			main_genericstandalone_rtio_core_sed_record104_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record88_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record88_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record88_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record88_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_address <= main_genericstandalone_rtio_core_sed_record88_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_data <= main_genericstandalone_rtio_core_sed_record88_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record96_rec_valid <= main_genericstandalone_rtio_core_sed_record88_rec_valid;
			main_genericstandalone_rtio_core_sed_record96_rec_seqn <= main_genericstandalone_rtio_core_sed_record88_rec_seqn;
			main_genericstandalone_rtio_core_sed_record96_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record88_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record96_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record88_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record88_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record88_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_address <= main_genericstandalone_rtio_core_sed_record88_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record96_rec_payload_data <= main_genericstandalone_rtio_core_sed_record88_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record104_rec_valid <= main_genericstandalone_rtio_core_sed_record80_rec_valid;
			main_genericstandalone_rtio_core_sed_record104_rec_seqn <= main_genericstandalone_rtio_core_sed_record80_rec_seqn;
			main_genericstandalone_rtio_core_sed_record104_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record80_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record80_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record80_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record80_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_address <= main_genericstandalone_rtio_core_sed_record80_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record104_rec_payload_data <= main_genericstandalone_rtio_core_sed_record80_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record81_rec_valid), main_genericstandalone_rtio_core_sed_record81_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record89_rec_valid), main_genericstandalone_rtio_core_sed_record89_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record81_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record81_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record89_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record89_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record81_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record89_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record81_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record81_rec_seqn < main_genericstandalone_rtio_core_sed_record89_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record97_rec_valid <= main_genericstandalone_rtio_core_sed_record89_rec_valid;
			main_genericstandalone_rtio_core_sed_record97_rec_seqn <= main_genericstandalone_rtio_core_sed_record89_rec_seqn;
			main_genericstandalone_rtio_core_sed_record97_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record89_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record97_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record89_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_address <= main_genericstandalone_rtio_core_sed_record89_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_data <= main_genericstandalone_rtio_core_sed_record89_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record105_rec_valid <= main_genericstandalone_rtio_core_sed_record81_rec_valid;
			main_genericstandalone_rtio_core_sed_record105_rec_seqn <= main_genericstandalone_rtio_core_sed_record81_rec_seqn;
			main_genericstandalone_rtio_core_sed_record105_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record81_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record81_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_address <= main_genericstandalone_rtio_core_sed_record81_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_data <= main_genericstandalone_rtio_core_sed_record81_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record97_rec_valid <= main_genericstandalone_rtio_core_sed_record81_rec_valid;
			main_genericstandalone_rtio_core_sed_record97_rec_seqn <= main_genericstandalone_rtio_core_sed_record81_rec_seqn;
			main_genericstandalone_rtio_core_sed_record97_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record81_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record97_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record81_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_address <= main_genericstandalone_rtio_core_sed_record81_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_data <= main_genericstandalone_rtio_core_sed_record81_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record105_rec_valid <= main_genericstandalone_rtio_core_sed_record89_rec_valid;
			main_genericstandalone_rtio_core_sed_record105_rec_seqn <= main_genericstandalone_rtio_core_sed_record89_rec_seqn;
			main_genericstandalone_rtio_core_sed_record105_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record89_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record89_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_address <= main_genericstandalone_rtio_core_sed_record89_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_data <= main_genericstandalone_rtio_core_sed_record89_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record97_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record97_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference39;
		main_genericstandalone_rtio_core_sed_record105_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record81_rec_valid), main_genericstandalone_rtio_core_sed_record81_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record89_rec_valid), main_genericstandalone_rtio_core_sed_record89_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record97_rec_valid <= main_genericstandalone_rtio_core_sed_record81_rec_valid;
			main_genericstandalone_rtio_core_sed_record97_rec_seqn <= main_genericstandalone_rtio_core_sed_record81_rec_seqn;
			main_genericstandalone_rtio_core_sed_record97_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record81_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record97_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record81_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_address <= main_genericstandalone_rtio_core_sed_record81_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_data <= main_genericstandalone_rtio_core_sed_record81_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record105_rec_valid <= main_genericstandalone_rtio_core_sed_record89_rec_valid;
			main_genericstandalone_rtio_core_sed_record105_rec_seqn <= main_genericstandalone_rtio_core_sed_record89_rec_seqn;
			main_genericstandalone_rtio_core_sed_record105_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record89_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record89_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_address <= main_genericstandalone_rtio_core_sed_record89_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_data <= main_genericstandalone_rtio_core_sed_record89_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record97_rec_valid <= main_genericstandalone_rtio_core_sed_record89_rec_valid;
			main_genericstandalone_rtio_core_sed_record97_rec_seqn <= main_genericstandalone_rtio_core_sed_record89_rec_seqn;
			main_genericstandalone_rtio_core_sed_record97_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record89_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record97_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record89_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record89_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record89_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_address <= main_genericstandalone_rtio_core_sed_record89_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record97_rec_payload_data <= main_genericstandalone_rtio_core_sed_record89_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record105_rec_valid <= main_genericstandalone_rtio_core_sed_record81_rec_valid;
			main_genericstandalone_rtio_core_sed_record105_rec_seqn <= main_genericstandalone_rtio_core_sed_record81_rec_seqn;
			main_genericstandalone_rtio_core_sed_record105_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record81_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record81_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record81_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record81_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_address <= main_genericstandalone_rtio_core_sed_record81_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record105_rec_payload_data <= main_genericstandalone_rtio_core_sed_record81_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record82_rec_valid), main_genericstandalone_rtio_core_sed_record82_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record90_rec_valid), main_genericstandalone_rtio_core_sed_record90_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record82_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record82_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record90_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record90_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record82_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record90_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record82_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record82_rec_seqn < main_genericstandalone_rtio_core_sed_record90_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record98_rec_valid <= main_genericstandalone_rtio_core_sed_record90_rec_valid;
			main_genericstandalone_rtio_core_sed_record98_rec_seqn <= main_genericstandalone_rtio_core_sed_record90_rec_seqn;
			main_genericstandalone_rtio_core_sed_record98_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record90_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record98_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record90_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_address <= main_genericstandalone_rtio_core_sed_record90_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_data <= main_genericstandalone_rtio_core_sed_record90_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record106_rec_valid <= main_genericstandalone_rtio_core_sed_record82_rec_valid;
			main_genericstandalone_rtio_core_sed_record106_rec_seqn <= main_genericstandalone_rtio_core_sed_record82_rec_seqn;
			main_genericstandalone_rtio_core_sed_record106_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record82_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record82_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_address <= main_genericstandalone_rtio_core_sed_record82_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_data <= main_genericstandalone_rtio_core_sed_record82_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record98_rec_valid <= main_genericstandalone_rtio_core_sed_record82_rec_valid;
			main_genericstandalone_rtio_core_sed_record98_rec_seqn <= main_genericstandalone_rtio_core_sed_record82_rec_seqn;
			main_genericstandalone_rtio_core_sed_record98_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record82_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record98_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record82_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_address <= main_genericstandalone_rtio_core_sed_record82_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_data <= main_genericstandalone_rtio_core_sed_record82_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record106_rec_valid <= main_genericstandalone_rtio_core_sed_record90_rec_valid;
			main_genericstandalone_rtio_core_sed_record106_rec_seqn <= main_genericstandalone_rtio_core_sed_record90_rec_seqn;
			main_genericstandalone_rtio_core_sed_record106_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record90_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record90_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_address <= main_genericstandalone_rtio_core_sed_record90_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_data <= main_genericstandalone_rtio_core_sed_record90_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record98_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record98_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference40;
		main_genericstandalone_rtio_core_sed_record106_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record82_rec_valid), main_genericstandalone_rtio_core_sed_record82_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record90_rec_valid), main_genericstandalone_rtio_core_sed_record90_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record98_rec_valid <= main_genericstandalone_rtio_core_sed_record82_rec_valid;
			main_genericstandalone_rtio_core_sed_record98_rec_seqn <= main_genericstandalone_rtio_core_sed_record82_rec_seqn;
			main_genericstandalone_rtio_core_sed_record98_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record82_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record98_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record82_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_address <= main_genericstandalone_rtio_core_sed_record82_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_data <= main_genericstandalone_rtio_core_sed_record82_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record106_rec_valid <= main_genericstandalone_rtio_core_sed_record90_rec_valid;
			main_genericstandalone_rtio_core_sed_record106_rec_seqn <= main_genericstandalone_rtio_core_sed_record90_rec_seqn;
			main_genericstandalone_rtio_core_sed_record106_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record90_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record90_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_address <= main_genericstandalone_rtio_core_sed_record90_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_data <= main_genericstandalone_rtio_core_sed_record90_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record98_rec_valid <= main_genericstandalone_rtio_core_sed_record90_rec_valid;
			main_genericstandalone_rtio_core_sed_record98_rec_seqn <= main_genericstandalone_rtio_core_sed_record90_rec_seqn;
			main_genericstandalone_rtio_core_sed_record98_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record90_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record98_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record90_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record90_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record90_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_address <= main_genericstandalone_rtio_core_sed_record90_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record98_rec_payload_data <= main_genericstandalone_rtio_core_sed_record90_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record106_rec_valid <= main_genericstandalone_rtio_core_sed_record82_rec_valid;
			main_genericstandalone_rtio_core_sed_record106_rec_seqn <= main_genericstandalone_rtio_core_sed_record82_rec_seqn;
			main_genericstandalone_rtio_core_sed_record106_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record82_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record82_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record82_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record82_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_address <= main_genericstandalone_rtio_core_sed_record82_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record106_rec_payload_data <= main_genericstandalone_rtio_core_sed_record82_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record83_rec_valid), main_genericstandalone_rtio_core_sed_record83_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record91_rec_valid), main_genericstandalone_rtio_core_sed_record91_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record83_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record83_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record91_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record91_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record83_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record91_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record83_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record83_rec_seqn < main_genericstandalone_rtio_core_sed_record91_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record99_rec_valid <= main_genericstandalone_rtio_core_sed_record91_rec_valid;
			main_genericstandalone_rtio_core_sed_record99_rec_seqn <= main_genericstandalone_rtio_core_sed_record91_rec_seqn;
			main_genericstandalone_rtio_core_sed_record99_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record91_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record99_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record91_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_address <= main_genericstandalone_rtio_core_sed_record91_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_data <= main_genericstandalone_rtio_core_sed_record91_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record107_rec_valid <= main_genericstandalone_rtio_core_sed_record83_rec_valid;
			main_genericstandalone_rtio_core_sed_record107_rec_seqn <= main_genericstandalone_rtio_core_sed_record83_rec_seqn;
			main_genericstandalone_rtio_core_sed_record107_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record83_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record83_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_address <= main_genericstandalone_rtio_core_sed_record83_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_data <= main_genericstandalone_rtio_core_sed_record83_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record99_rec_valid <= main_genericstandalone_rtio_core_sed_record83_rec_valid;
			main_genericstandalone_rtio_core_sed_record99_rec_seqn <= main_genericstandalone_rtio_core_sed_record83_rec_seqn;
			main_genericstandalone_rtio_core_sed_record99_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record83_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record99_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record83_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_address <= main_genericstandalone_rtio_core_sed_record83_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_data <= main_genericstandalone_rtio_core_sed_record83_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record107_rec_valid <= main_genericstandalone_rtio_core_sed_record91_rec_valid;
			main_genericstandalone_rtio_core_sed_record107_rec_seqn <= main_genericstandalone_rtio_core_sed_record91_rec_seqn;
			main_genericstandalone_rtio_core_sed_record107_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record91_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record91_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_address <= main_genericstandalone_rtio_core_sed_record91_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_data <= main_genericstandalone_rtio_core_sed_record91_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record99_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record99_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference41;
		main_genericstandalone_rtio_core_sed_record107_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record83_rec_valid), main_genericstandalone_rtio_core_sed_record83_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record91_rec_valid), main_genericstandalone_rtio_core_sed_record91_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record99_rec_valid <= main_genericstandalone_rtio_core_sed_record83_rec_valid;
			main_genericstandalone_rtio_core_sed_record99_rec_seqn <= main_genericstandalone_rtio_core_sed_record83_rec_seqn;
			main_genericstandalone_rtio_core_sed_record99_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record83_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record99_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record83_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_address <= main_genericstandalone_rtio_core_sed_record83_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_data <= main_genericstandalone_rtio_core_sed_record83_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record107_rec_valid <= main_genericstandalone_rtio_core_sed_record91_rec_valid;
			main_genericstandalone_rtio_core_sed_record107_rec_seqn <= main_genericstandalone_rtio_core_sed_record91_rec_seqn;
			main_genericstandalone_rtio_core_sed_record107_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record91_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record91_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_address <= main_genericstandalone_rtio_core_sed_record91_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_data <= main_genericstandalone_rtio_core_sed_record91_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record99_rec_valid <= main_genericstandalone_rtio_core_sed_record91_rec_valid;
			main_genericstandalone_rtio_core_sed_record99_rec_seqn <= main_genericstandalone_rtio_core_sed_record91_rec_seqn;
			main_genericstandalone_rtio_core_sed_record99_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record91_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record99_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record91_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record91_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record91_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_address <= main_genericstandalone_rtio_core_sed_record91_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record99_rec_payload_data <= main_genericstandalone_rtio_core_sed_record91_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record107_rec_valid <= main_genericstandalone_rtio_core_sed_record83_rec_valid;
			main_genericstandalone_rtio_core_sed_record107_rec_seqn <= main_genericstandalone_rtio_core_sed_record83_rec_seqn;
			main_genericstandalone_rtio_core_sed_record107_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record83_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record83_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record83_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record83_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_address <= main_genericstandalone_rtio_core_sed_record83_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record107_rec_payload_data <= main_genericstandalone_rtio_core_sed_record83_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record84_rec_valid), main_genericstandalone_rtio_core_sed_record84_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record92_rec_valid), main_genericstandalone_rtio_core_sed_record92_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record84_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record84_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record92_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record92_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record84_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record92_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record84_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record84_rec_seqn < main_genericstandalone_rtio_core_sed_record92_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record100_rec_valid <= main_genericstandalone_rtio_core_sed_record92_rec_valid;
			main_genericstandalone_rtio_core_sed_record100_rec_seqn <= main_genericstandalone_rtio_core_sed_record92_rec_seqn;
			main_genericstandalone_rtio_core_sed_record100_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record92_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record92_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_address <= main_genericstandalone_rtio_core_sed_record92_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_data <= main_genericstandalone_rtio_core_sed_record92_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record108_rec_valid <= main_genericstandalone_rtio_core_sed_record84_rec_valid;
			main_genericstandalone_rtio_core_sed_record108_rec_seqn <= main_genericstandalone_rtio_core_sed_record84_rec_seqn;
			main_genericstandalone_rtio_core_sed_record108_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record84_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record108_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record84_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_address <= main_genericstandalone_rtio_core_sed_record84_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_data <= main_genericstandalone_rtio_core_sed_record84_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record100_rec_valid <= main_genericstandalone_rtio_core_sed_record84_rec_valid;
			main_genericstandalone_rtio_core_sed_record100_rec_seqn <= main_genericstandalone_rtio_core_sed_record84_rec_seqn;
			main_genericstandalone_rtio_core_sed_record100_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record84_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record84_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_address <= main_genericstandalone_rtio_core_sed_record84_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_data <= main_genericstandalone_rtio_core_sed_record84_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record108_rec_valid <= main_genericstandalone_rtio_core_sed_record92_rec_valid;
			main_genericstandalone_rtio_core_sed_record108_rec_seqn <= main_genericstandalone_rtio_core_sed_record92_rec_seqn;
			main_genericstandalone_rtio_core_sed_record108_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record92_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record108_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record92_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_address <= main_genericstandalone_rtio_core_sed_record92_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_data <= main_genericstandalone_rtio_core_sed_record92_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record100_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference42;
		main_genericstandalone_rtio_core_sed_record108_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record84_rec_valid), main_genericstandalone_rtio_core_sed_record84_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record92_rec_valid), main_genericstandalone_rtio_core_sed_record92_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record100_rec_valid <= main_genericstandalone_rtio_core_sed_record84_rec_valid;
			main_genericstandalone_rtio_core_sed_record100_rec_seqn <= main_genericstandalone_rtio_core_sed_record84_rec_seqn;
			main_genericstandalone_rtio_core_sed_record100_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record84_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record84_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_address <= main_genericstandalone_rtio_core_sed_record84_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_data <= main_genericstandalone_rtio_core_sed_record84_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record108_rec_valid <= main_genericstandalone_rtio_core_sed_record92_rec_valid;
			main_genericstandalone_rtio_core_sed_record108_rec_seqn <= main_genericstandalone_rtio_core_sed_record92_rec_seqn;
			main_genericstandalone_rtio_core_sed_record108_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record92_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record108_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record92_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_address <= main_genericstandalone_rtio_core_sed_record92_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_data <= main_genericstandalone_rtio_core_sed_record92_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record100_rec_valid <= main_genericstandalone_rtio_core_sed_record92_rec_valid;
			main_genericstandalone_rtio_core_sed_record100_rec_seqn <= main_genericstandalone_rtio_core_sed_record92_rec_seqn;
			main_genericstandalone_rtio_core_sed_record100_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record92_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record92_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record92_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record92_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_address <= main_genericstandalone_rtio_core_sed_record92_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record100_rec_payload_data <= main_genericstandalone_rtio_core_sed_record92_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record108_rec_valid <= main_genericstandalone_rtio_core_sed_record84_rec_valid;
			main_genericstandalone_rtio_core_sed_record108_rec_seqn <= main_genericstandalone_rtio_core_sed_record84_rec_seqn;
			main_genericstandalone_rtio_core_sed_record108_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record84_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record108_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record84_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record84_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record84_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_address <= main_genericstandalone_rtio_core_sed_record84_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record108_rec_payload_data <= main_genericstandalone_rtio_core_sed_record84_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record85_rec_valid), main_genericstandalone_rtio_core_sed_record85_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record93_rec_valid), main_genericstandalone_rtio_core_sed_record93_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record85_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record85_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record93_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record93_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record85_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record93_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record85_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record85_rec_seqn < main_genericstandalone_rtio_core_sed_record93_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record101_rec_valid <= main_genericstandalone_rtio_core_sed_record93_rec_valid;
			main_genericstandalone_rtio_core_sed_record101_rec_seqn <= main_genericstandalone_rtio_core_sed_record93_rec_seqn;
			main_genericstandalone_rtio_core_sed_record101_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record93_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record93_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_address <= main_genericstandalone_rtio_core_sed_record93_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_data <= main_genericstandalone_rtio_core_sed_record93_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record109_rec_valid <= main_genericstandalone_rtio_core_sed_record85_rec_valid;
			main_genericstandalone_rtio_core_sed_record109_rec_seqn <= main_genericstandalone_rtio_core_sed_record85_rec_seqn;
			main_genericstandalone_rtio_core_sed_record109_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record85_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record109_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record85_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_address <= main_genericstandalone_rtio_core_sed_record85_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_data <= main_genericstandalone_rtio_core_sed_record85_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record101_rec_valid <= main_genericstandalone_rtio_core_sed_record85_rec_valid;
			main_genericstandalone_rtio_core_sed_record101_rec_seqn <= main_genericstandalone_rtio_core_sed_record85_rec_seqn;
			main_genericstandalone_rtio_core_sed_record101_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record85_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record85_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_address <= main_genericstandalone_rtio_core_sed_record85_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_data <= main_genericstandalone_rtio_core_sed_record85_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record109_rec_valid <= main_genericstandalone_rtio_core_sed_record93_rec_valid;
			main_genericstandalone_rtio_core_sed_record109_rec_seqn <= main_genericstandalone_rtio_core_sed_record93_rec_seqn;
			main_genericstandalone_rtio_core_sed_record109_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record93_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record109_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record93_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_address <= main_genericstandalone_rtio_core_sed_record93_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_data <= main_genericstandalone_rtio_core_sed_record93_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record101_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference43;
		main_genericstandalone_rtio_core_sed_record109_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record85_rec_valid), main_genericstandalone_rtio_core_sed_record85_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record93_rec_valid), main_genericstandalone_rtio_core_sed_record93_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record101_rec_valid <= main_genericstandalone_rtio_core_sed_record85_rec_valid;
			main_genericstandalone_rtio_core_sed_record101_rec_seqn <= main_genericstandalone_rtio_core_sed_record85_rec_seqn;
			main_genericstandalone_rtio_core_sed_record101_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record85_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record85_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_address <= main_genericstandalone_rtio_core_sed_record85_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_data <= main_genericstandalone_rtio_core_sed_record85_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record109_rec_valid <= main_genericstandalone_rtio_core_sed_record93_rec_valid;
			main_genericstandalone_rtio_core_sed_record109_rec_seqn <= main_genericstandalone_rtio_core_sed_record93_rec_seqn;
			main_genericstandalone_rtio_core_sed_record109_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record93_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record109_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record93_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_address <= main_genericstandalone_rtio_core_sed_record93_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_data <= main_genericstandalone_rtio_core_sed_record93_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record101_rec_valid <= main_genericstandalone_rtio_core_sed_record93_rec_valid;
			main_genericstandalone_rtio_core_sed_record101_rec_seqn <= main_genericstandalone_rtio_core_sed_record93_rec_seqn;
			main_genericstandalone_rtio_core_sed_record101_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record93_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record93_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record93_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record93_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_address <= main_genericstandalone_rtio_core_sed_record93_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record101_rec_payload_data <= main_genericstandalone_rtio_core_sed_record93_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record109_rec_valid <= main_genericstandalone_rtio_core_sed_record85_rec_valid;
			main_genericstandalone_rtio_core_sed_record109_rec_seqn <= main_genericstandalone_rtio_core_sed_record85_rec_seqn;
			main_genericstandalone_rtio_core_sed_record109_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record85_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record109_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record85_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record85_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record85_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_address <= main_genericstandalone_rtio_core_sed_record85_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record109_rec_payload_data <= main_genericstandalone_rtio_core_sed_record85_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record86_rec_valid), main_genericstandalone_rtio_core_sed_record86_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record94_rec_valid), main_genericstandalone_rtio_core_sed_record94_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record86_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record86_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record94_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record94_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record86_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record94_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record86_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record86_rec_seqn < main_genericstandalone_rtio_core_sed_record94_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record102_rec_valid <= main_genericstandalone_rtio_core_sed_record94_rec_valid;
			main_genericstandalone_rtio_core_sed_record102_rec_seqn <= main_genericstandalone_rtio_core_sed_record94_rec_seqn;
			main_genericstandalone_rtio_core_sed_record102_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record94_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record94_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_address <= main_genericstandalone_rtio_core_sed_record94_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_data <= main_genericstandalone_rtio_core_sed_record94_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record110_rec_valid <= main_genericstandalone_rtio_core_sed_record86_rec_valid;
			main_genericstandalone_rtio_core_sed_record110_rec_seqn <= main_genericstandalone_rtio_core_sed_record86_rec_seqn;
			main_genericstandalone_rtio_core_sed_record110_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record86_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record110_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record86_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_address <= main_genericstandalone_rtio_core_sed_record86_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_data <= main_genericstandalone_rtio_core_sed_record86_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record102_rec_valid <= main_genericstandalone_rtio_core_sed_record86_rec_valid;
			main_genericstandalone_rtio_core_sed_record102_rec_seqn <= main_genericstandalone_rtio_core_sed_record86_rec_seqn;
			main_genericstandalone_rtio_core_sed_record102_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record86_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record86_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_address <= main_genericstandalone_rtio_core_sed_record86_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_data <= main_genericstandalone_rtio_core_sed_record86_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record110_rec_valid <= main_genericstandalone_rtio_core_sed_record94_rec_valid;
			main_genericstandalone_rtio_core_sed_record110_rec_seqn <= main_genericstandalone_rtio_core_sed_record94_rec_seqn;
			main_genericstandalone_rtio_core_sed_record110_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record94_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record110_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record94_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_address <= main_genericstandalone_rtio_core_sed_record94_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_data <= main_genericstandalone_rtio_core_sed_record94_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record102_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference44;
		main_genericstandalone_rtio_core_sed_record110_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record86_rec_valid), main_genericstandalone_rtio_core_sed_record86_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record94_rec_valid), main_genericstandalone_rtio_core_sed_record94_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record102_rec_valid <= main_genericstandalone_rtio_core_sed_record86_rec_valid;
			main_genericstandalone_rtio_core_sed_record102_rec_seqn <= main_genericstandalone_rtio_core_sed_record86_rec_seqn;
			main_genericstandalone_rtio_core_sed_record102_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record86_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record86_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_address <= main_genericstandalone_rtio_core_sed_record86_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_data <= main_genericstandalone_rtio_core_sed_record86_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record110_rec_valid <= main_genericstandalone_rtio_core_sed_record94_rec_valid;
			main_genericstandalone_rtio_core_sed_record110_rec_seqn <= main_genericstandalone_rtio_core_sed_record94_rec_seqn;
			main_genericstandalone_rtio_core_sed_record110_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record94_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record110_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record94_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_address <= main_genericstandalone_rtio_core_sed_record94_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_data <= main_genericstandalone_rtio_core_sed_record94_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record102_rec_valid <= main_genericstandalone_rtio_core_sed_record94_rec_valid;
			main_genericstandalone_rtio_core_sed_record102_rec_seqn <= main_genericstandalone_rtio_core_sed_record94_rec_seqn;
			main_genericstandalone_rtio_core_sed_record102_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record94_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record94_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record94_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record94_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_address <= main_genericstandalone_rtio_core_sed_record94_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record102_rec_payload_data <= main_genericstandalone_rtio_core_sed_record94_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record110_rec_valid <= main_genericstandalone_rtio_core_sed_record86_rec_valid;
			main_genericstandalone_rtio_core_sed_record110_rec_seqn <= main_genericstandalone_rtio_core_sed_record86_rec_seqn;
			main_genericstandalone_rtio_core_sed_record110_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record86_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record110_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record86_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record86_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record86_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_address <= main_genericstandalone_rtio_core_sed_record86_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record110_rec_payload_data <= main_genericstandalone_rtio_core_sed_record86_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record87_rec_valid), main_genericstandalone_rtio_core_sed_record87_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record95_rec_valid), main_genericstandalone_rtio_core_sed_record95_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record87_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record87_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record95_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record95_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record87_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record95_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record87_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record87_rec_seqn < main_genericstandalone_rtio_core_sed_record95_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record103_rec_valid <= main_genericstandalone_rtio_core_sed_record95_rec_valid;
			main_genericstandalone_rtio_core_sed_record103_rec_seqn <= main_genericstandalone_rtio_core_sed_record95_rec_seqn;
			main_genericstandalone_rtio_core_sed_record103_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record95_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record95_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record95_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record95_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_address <= main_genericstandalone_rtio_core_sed_record95_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_data <= main_genericstandalone_rtio_core_sed_record95_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record111_rec_valid <= main_genericstandalone_rtio_core_sed_record87_rec_valid;
			main_genericstandalone_rtio_core_sed_record111_rec_seqn <= main_genericstandalone_rtio_core_sed_record87_rec_seqn;
			main_genericstandalone_rtio_core_sed_record111_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record87_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record111_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record87_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record87_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record87_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_address <= main_genericstandalone_rtio_core_sed_record87_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_data <= main_genericstandalone_rtio_core_sed_record87_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record103_rec_valid <= main_genericstandalone_rtio_core_sed_record87_rec_valid;
			main_genericstandalone_rtio_core_sed_record103_rec_seqn <= main_genericstandalone_rtio_core_sed_record87_rec_seqn;
			main_genericstandalone_rtio_core_sed_record103_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record87_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record87_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record87_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record87_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_address <= main_genericstandalone_rtio_core_sed_record87_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_data <= main_genericstandalone_rtio_core_sed_record87_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record111_rec_valid <= main_genericstandalone_rtio_core_sed_record95_rec_valid;
			main_genericstandalone_rtio_core_sed_record111_rec_seqn <= main_genericstandalone_rtio_core_sed_record95_rec_seqn;
			main_genericstandalone_rtio_core_sed_record111_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record95_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record111_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record95_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record95_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record95_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_address <= main_genericstandalone_rtio_core_sed_record95_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_data <= main_genericstandalone_rtio_core_sed_record95_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record103_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference45;
		main_genericstandalone_rtio_core_sed_record111_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record87_rec_valid), main_genericstandalone_rtio_core_sed_record87_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record95_rec_valid), main_genericstandalone_rtio_core_sed_record95_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record103_rec_valid <= main_genericstandalone_rtio_core_sed_record87_rec_valid;
			main_genericstandalone_rtio_core_sed_record103_rec_seqn <= main_genericstandalone_rtio_core_sed_record87_rec_seqn;
			main_genericstandalone_rtio_core_sed_record103_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record87_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record87_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record87_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record87_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_address <= main_genericstandalone_rtio_core_sed_record87_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_data <= main_genericstandalone_rtio_core_sed_record87_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record111_rec_valid <= main_genericstandalone_rtio_core_sed_record95_rec_valid;
			main_genericstandalone_rtio_core_sed_record111_rec_seqn <= main_genericstandalone_rtio_core_sed_record95_rec_seqn;
			main_genericstandalone_rtio_core_sed_record111_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record95_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record111_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record95_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record95_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record95_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_address <= main_genericstandalone_rtio_core_sed_record95_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_data <= main_genericstandalone_rtio_core_sed_record95_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record103_rec_valid <= main_genericstandalone_rtio_core_sed_record95_rec_valid;
			main_genericstandalone_rtio_core_sed_record103_rec_seqn <= main_genericstandalone_rtio_core_sed_record95_rec_seqn;
			main_genericstandalone_rtio_core_sed_record103_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record95_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record95_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record95_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record95_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_address <= main_genericstandalone_rtio_core_sed_record95_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record103_rec_payload_data <= main_genericstandalone_rtio_core_sed_record95_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record111_rec_valid <= main_genericstandalone_rtio_core_sed_record87_rec_valid;
			main_genericstandalone_rtio_core_sed_record111_rec_seqn <= main_genericstandalone_rtio_core_sed_record87_rec_seqn;
			main_genericstandalone_rtio_core_sed_record111_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record87_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record111_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record87_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record87_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record87_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_address <= main_genericstandalone_rtio_core_sed_record87_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record111_rec_payload_data <= main_genericstandalone_rtio_core_sed_record87_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record100_rec_valid), main_genericstandalone_rtio_core_sed_record100_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record104_rec_valid), main_genericstandalone_rtio_core_sed_record104_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record100_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record100_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record104_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record104_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record100_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record104_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record100_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record100_rec_seqn < main_genericstandalone_rtio_core_sed_record104_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record116_rec_valid <= main_genericstandalone_rtio_core_sed_record104_rec_valid;
			main_genericstandalone_rtio_core_sed_record116_rec_seqn <= main_genericstandalone_rtio_core_sed_record104_rec_seqn;
			main_genericstandalone_rtio_core_sed_record116_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record104_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record104_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_address <= main_genericstandalone_rtio_core_sed_record104_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_data <= main_genericstandalone_rtio_core_sed_record104_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record120_rec_valid <= main_genericstandalone_rtio_core_sed_record100_rec_valid;
			main_genericstandalone_rtio_core_sed_record120_rec_seqn <= main_genericstandalone_rtio_core_sed_record100_rec_seqn;
			main_genericstandalone_rtio_core_sed_record120_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record100_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record100_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_address <= main_genericstandalone_rtio_core_sed_record100_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_data <= main_genericstandalone_rtio_core_sed_record100_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record116_rec_valid <= main_genericstandalone_rtio_core_sed_record100_rec_valid;
			main_genericstandalone_rtio_core_sed_record116_rec_seqn <= main_genericstandalone_rtio_core_sed_record100_rec_seqn;
			main_genericstandalone_rtio_core_sed_record116_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record100_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record100_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_address <= main_genericstandalone_rtio_core_sed_record100_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_data <= main_genericstandalone_rtio_core_sed_record100_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record120_rec_valid <= main_genericstandalone_rtio_core_sed_record104_rec_valid;
			main_genericstandalone_rtio_core_sed_record120_rec_seqn <= main_genericstandalone_rtio_core_sed_record104_rec_seqn;
			main_genericstandalone_rtio_core_sed_record120_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record104_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record104_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_address <= main_genericstandalone_rtio_core_sed_record104_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_data <= main_genericstandalone_rtio_core_sed_record104_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record116_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference46;
		main_genericstandalone_rtio_core_sed_record120_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record100_rec_valid), main_genericstandalone_rtio_core_sed_record100_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record104_rec_valid), main_genericstandalone_rtio_core_sed_record104_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record116_rec_valid <= main_genericstandalone_rtio_core_sed_record100_rec_valid;
			main_genericstandalone_rtio_core_sed_record116_rec_seqn <= main_genericstandalone_rtio_core_sed_record100_rec_seqn;
			main_genericstandalone_rtio_core_sed_record116_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record100_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record100_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_address <= main_genericstandalone_rtio_core_sed_record100_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_data <= main_genericstandalone_rtio_core_sed_record100_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record120_rec_valid <= main_genericstandalone_rtio_core_sed_record104_rec_valid;
			main_genericstandalone_rtio_core_sed_record120_rec_seqn <= main_genericstandalone_rtio_core_sed_record104_rec_seqn;
			main_genericstandalone_rtio_core_sed_record120_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record104_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record104_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_address <= main_genericstandalone_rtio_core_sed_record104_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_data <= main_genericstandalone_rtio_core_sed_record104_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record116_rec_valid <= main_genericstandalone_rtio_core_sed_record104_rec_valid;
			main_genericstandalone_rtio_core_sed_record116_rec_seqn <= main_genericstandalone_rtio_core_sed_record104_rec_seqn;
			main_genericstandalone_rtio_core_sed_record116_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record104_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record104_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record104_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record104_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_address <= main_genericstandalone_rtio_core_sed_record104_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record116_rec_payload_data <= main_genericstandalone_rtio_core_sed_record104_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record120_rec_valid <= main_genericstandalone_rtio_core_sed_record100_rec_valid;
			main_genericstandalone_rtio_core_sed_record120_rec_seqn <= main_genericstandalone_rtio_core_sed_record100_rec_seqn;
			main_genericstandalone_rtio_core_sed_record120_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record100_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record100_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record100_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record100_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_address <= main_genericstandalone_rtio_core_sed_record100_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record120_rec_payload_data <= main_genericstandalone_rtio_core_sed_record100_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record101_rec_valid), main_genericstandalone_rtio_core_sed_record101_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record105_rec_valid), main_genericstandalone_rtio_core_sed_record105_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record101_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record101_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record105_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record105_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record101_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record105_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record101_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record101_rec_seqn < main_genericstandalone_rtio_core_sed_record105_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record117_rec_valid <= main_genericstandalone_rtio_core_sed_record105_rec_valid;
			main_genericstandalone_rtio_core_sed_record117_rec_seqn <= main_genericstandalone_rtio_core_sed_record105_rec_seqn;
			main_genericstandalone_rtio_core_sed_record117_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record105_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record105_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_address <= main_genericstandalone_rtio_core_sed_record105_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_data <= main_genericstandalone_rtio_core_sed_record105_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record121_rec_valid <= main_genericstandalone_rtio_core_sed_record101_rec_valid;
			main_genericstandalone_rtio_core_sed_record121_rec_seqn <= main_genericstandalone_rtio_core_sed_record101_rec_seqn;
			main_genericstandalone_rtio_core_sed_record121_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record101_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record101_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_address <= main_genericstandalone_rtio_core_sed_record101_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_data <= main_genericstandalone_rtio_core_sed_record101_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record117_rec_valid <= main_genericstandalone_rtio_core_sed_record101_rec_valid;
			main_genericstandalone_rtio_core_sed_record117_rec_seqn <= main_genericstandalone_rtio_core_sed_record101_rec_seqn;
			main_genericstandalone_rtio_core_sed_record117_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record101_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record101_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_address <= main_genericstandalone_rtio_core_sed_record101_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_data <= main_genericstandalone_rtio_core_sed_record101_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record121_rec_valid <= main_genericstandalone_rtio_core_sed_record105_rec_valid;
			main_genericstandalone_rtio_core_sed_record121_rec_seqn <= main_genericstandalone_rtio_core_sed_record105_rec_seqn;
			main_genericstandalone_rtio_core_sed_record121_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record105_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record105_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_address <= main_genericstandalone_rtio_core_sed_record105_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_data <= main_genericstandalone_rtio_core_sed_record105_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record117_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference47;
		main_genericstandalone_rtio_core_sed_record121_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record101_rec_valid), main_genericstandalone_rtio_core_sed_record101_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record105_rec_valid), main_genericstandalone_rtio_core_sed_record105_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record117_rec_valid <= main_genericstandalone_rtio_core_sed_record101_rec_valid;
			main_genericstandalone_rtio_core_sed_record117_rec_seqn <= main_genericstandalone_rtio_core_sed_record101_rec_seqn;
			main_genericstandalone_rtio_core_sed_record117_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record101_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record101_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_address <= main_genericstandalone_rtio_core_sed_record101_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_data <= main_genericstandalone_rtio_core_sed_record101_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record121_rec_valid <= main_genericstandalone_rtio_core_sed_record105_rec_valid;
			main_genericstandalone_rtio_core_sed_record121_rec_seqn <= main_genericstandalone_rtio_core_sed_record105_rec_seqn;
			main_genericstandalone_rtio_core_sed_record121_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record105_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record105_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_address <= main_genericstandalone_rtio_core_sed_record105_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_data <= main_genericstandalone_rtio_core_sed_record105_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record117_rec_valid <= main_genericstandalone_rtio_core_sed_record105_rec_valid;
			main_genericstandalone_rtio_core_sed_record117_rec_seqn <= main_genericstandalone_rtio_core_sed_record105_rec_seqn;
			main_genericstandalone_rtio_core_sed_record117_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record105_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record105_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record105_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record105_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_address <= main_genericstandalone_rtio_core_sed_record105_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record117_rec_payload_data <= main_genericstandalone_rtio_core_sed_record105_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record121_rec_valid <= main_genericstandalone_rtio_core_sed_record101_rec_valid;
			main_genericstandalone_rtio_core_sed_record121_rec_seqn <= main_genericstandalone_rtio_core_sed_record101_rec_seqn;
			main_genericstandalone_rtio_core_sed_record121_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record101_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record101_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record101_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record101_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_address <= main_genericstandalone_rtio_core_sed_record101_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record121_rec_payload_data <= main_genericstandalone_rtio_core_sed_record101_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record102_rec_valid), main_genericstandalone_rtio_core_sed_record102_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record106_rec_valid), main_genericstandalone_rtio_core_sed_record106_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record102_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record102_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record106_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record106_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record102_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record106_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record102_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record102_rec_seqn < main_genericstandalone_rtio_core_sed_record106_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record118_rec_valid <= main_genericstandalone_rtio_core_sed_record106_rec_valid;
			main_genericstandalone_rtio_core_sed_record118_rec_seqn <= main_genericstandalone_rtio_core_sed_record106_rec_seqn;
			main_genericstandalone_rtio_core_sed_record118_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record106_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record106_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_address <= main_genericstandalone_rtio_core_sed_record106_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_data <= main_genericstandalone_rtio_core_sed_record106_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record122_rec_valid <= main_genericstandalone_rtio_core_sed_record102_rec_valid;
			main_genericstandalone_rtio_core_sed_record122_rec_seqn <= main_genericstandalone_rtio_core_sed_record102_rec_seqn;
			main_genericstandalone_rtio_core_sed_record122_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record102_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record102_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_address <= main_genericstandalone_rtio_core_sed_record102_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_data <= main_genericstandalone_rtio_core_sed_record102_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record118_rec_valid <= main_genericstandalone_rtio_core_sed_record102_rec_valid;
			main_genericstandalone_rtio_core_sed_record118_rec_seqn <= main_genericstandalone_rtio_core_sed_record102_rec_seqn;
			main_genericstandalone_rtio_core_sed_record118_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record102_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record102_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_address <= main_genericstandalone_rtio_core_sed_record102_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_data <= main_genericstandalone_rtio_core_sed_record102_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record122_rec_valid <= main_genericstandalone_rtio_core_sed_record106_rec_valid;
			main_genericstandalone_rtio_core_sed_record122_rec_seqn <= main_genericstandalone_rtio_core_sed_record106_rec_seqn;
			main_genericstandalone_rtio_core_sed_record122_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record106_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record106_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_address <= main_genericstandalone_rtio_core_sed_record106_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_data <= main_genericstandalone_rtio_core_sed_record106_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record118_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference48;
		main_genericstandalone_rtio_core_sed_record122_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record102_rec_valid), main_genericstandalone_rtio_core_sed_record102_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record106_rec_valid), main_genericstandalone_rtio_core_sed_record106_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record118_rec_valid <= main_genericstandalone_rtio_core_sed_record102_rec_valid;
			main_genericstandalone_rtio_core_sed_record118_rec_seqn <= main_genericstandalone_rtio_core_sed_record102_rec_seqn;
			main_genericstandalone_rtio_core_sed_record118_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record102_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record102_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_address <= main_genericstandalone_rtio_core_sed_record102_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_data <= main_genericstandalone_rtio_core_sed_record102_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record122_rec_valid <= main_genericstandalone_rtio_core_sed_record106_rec_valid;
			main_genericstandalone_rtio_core_sed_record122_rec_seqn <= main_genericstandalone_rtio_core_sed_record106_rec_seqn;
			main_genericstandalone_rtio_core_sed_record122_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record106_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record106_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_address <= main_genericstandalone_rtio_core_sed_record106_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_data <= main_genericstandalone_rtio_core_sed_record106_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record118_rec_valid <= main_genericstandalone_rtio_core_sed_record106_rec_valid;
			main_genericstandalone_rtio_core_sed_record118_rec_seqn <= main_genericstandalone_rtio_core_sed_record106_rec_seqn;
			main_genericstandalone_rtio_core_sed_record118_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record106_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record106_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record106_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record106_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_address <= main_genericstandalone_rtio_core_sed_record106_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record118_rec_payload_data <= main_genericstandalone_rtio_core_sed_record106_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record122_rec_valid <= main_genericstandalone_rtio_core_sed_record102_rec_valid;
			main_genericstandalone_rtio_core_sed_record122_rec_seqn <= main_genericstandalone_rtio_core_sed_record102_rec_seqn;
			main_genericstandalone_rtio_core_sed_record122_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record102_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record102_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record102_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record102_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_address <= main_genericstandalone_rtio_core_sed_record102_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record122_rec_payload_data <= main_genericstandalone_rtio_core_sed_record102_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record103_rec_valid), main_genericstandalone_rtio_core_sed_record103_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record107_rec_valid), main_genericstandalone_rtio_core_sed_record107_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record103_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record103_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record107_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record107_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record103_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record107_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record103_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record103_rec_seqn < main_genericstandalone_rtio_core_sed_record107_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record119_rec_valid <= main_genericstandalone_rtio_core_sed_record107_rec_valid;
			main_genericstandalone_rtio_core_sed_record119_rec_seqn <= main_genericstandalone_rtio_core_sed_record107_rec_seqn;
			main_genericstandalone_rtio_core_sed_record119_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record107_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record107_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_address <= main_genericstandalone_rtio_core_sed_record107_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_data <= main_genericstandalone_rtio_core_sed_record107_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record123_rec_valid <= main_genericstandalone_rtio_core_sed_record103_rec_valid;
			main_genericstandalone_rtio_core_sed_record123_rec_seqn <= main_genericstandalone_rtio_core_sed_record103_rec_seqn;
			main_genericstandalone_rtio_core_sed_record123_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record103_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record103_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_address <= main_genericstandalone_rtio_core_sed_record103_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_data <= main_genericstandalone_rtio_core_sed_record103_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record119_rec_valid <= main_genericstandalone_rtio_core_sed_record103_rec_valid;
			main_genericstandalone_rtio_core_sed_record119_rec_seqn <= main_genericstandalone_rtio_core_sed_record103_rec_seqn;
			main_genericstandalone_rtio_core_sed_record119_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record103_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record103_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_address <= main_genericstandalone_rtio_core_sed_record103_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_data <= main_genericstandalone_rtio_core_sed_record103_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record123_rec_valid <= main_genericstandalone_rtio_core_sed_record107_rec_valid;
			main_genericstandalone_rtio_core_sed_record123_rec_seqn <= main_genericstandalone_rtio_core_sed_record107_rec_seqn;
			main_genericstandalone_rtio_core_sed_record123_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record107_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record107_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_address <= main_genericstandalone_rtio_core_sed_record107_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_data <= main_genericstandalone_rtio_core_sed_record107_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record119_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference49;
		main_genericstandalone_rtio_core_sed_record123_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record103_rec_valid), main_genericstandalone_rtio_core_sed_record103_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record107_rec_valid), main_genericstandalone_rtio_core_sed_record107_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record119_rec_valid <= main_genericstandalone_rtio_core_sed_record103_rec_valid;
			main_genericstandalone_rtio_core_sed_record119_rec_seqn <= main_genericstandalone_rtio_core_sed_record103_rec_seqn;
			main_genericstandalone_rtio_core_sed_record119_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record103_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record103_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_address <= main_genericstandalone_rtio_core_sed_record103_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_data <= main_genericstandalone_rtio_core_sed_record103_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record123_rec_valid <= main_genericstandalone_rtio_core_sed_record107_rec_valid;
			main_genericstandalone_rtio_core_sed_record123_rec_seqn <= main_genericstandalone_rtio_core_sed_record107_rec_seqn;
			main_genericstandalone_rtio_core_sed_record123_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record107_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record107_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_address <= main_genericstandalone_rtio_core_sed_record107_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_data <= main_genericstandalone_rtio_core_sed_record107_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record119_rec_valid <= main_genericstandalone_rtio_core_sed_record107_rec_valid;
			main_genericstandalone_rtio_core_sed_record119_rec_seqn <= main_genericstandalone_rtio_core_sed_record107_rec_seqn;
			main_genericstandalone_rtio_core_sed_record119_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record107_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record107_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record107_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record107_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_address <= main_genericstandalone_rtio_core_sed_record107_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record119_rec_payload_data <= main_genericstandalone_rtio_core_sed_record107_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record123_rec_valid <= main_genericstandalone_rtio_core_sed_record103_rec_valid;
			main_genericstandalone_rtio_core_sed_record123_rec_seqn <= main_genericstandalone_rtio_core_sed_record103_rec_seqn;
			main_genericstandalone_rtio_core_sed_record123_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record103_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record103_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record103_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record103_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_address <= main_genericstandalone_rtio_core_sed_record103_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record123_rec_payload_data <= main_genericstandalone_rtio_core_sed_record103_rec_payload_data;
		end
	end
	main_genericstandalone_rtio_core_sed_record112_rec_valid <= main_genericstandalone_rtio_core_sed_record96_rec_valid;
	main_genericstandalone_rtio_core_sed_record112_rec_seqn <= main_genericstandalone_rtio_core_sed_record96_rec_seqn;
	main_genericstandalone_rtio_core_sed_record112_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record96_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record112_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record96_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record112_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record96_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record112_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record96_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record112_rec_payload_address <= main_genericstandalone_rtio_core_sed_record96_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record112_rec_payload_data <= main_genericstandalone_rtio_core_sed_record96_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record113_rec_valid <= main_genericstandalone_rtio_core_sed_record97_rec_valid;
	main_genericstandalone_rtio_core_sed_record113_rec_seqn <= main_genericstandalone_rtio_core_sed_record97_rec_seqn;
	main_genericstandalone_rtio_core_sed_record113_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record97_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record113_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record97_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record113_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record97_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record113_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record97_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record113_rec_payload_address <= main_genericstandalone_rtio_core_sed_record97_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record113_rec_payload_data <= main_genericstandalone_rtio_core_sed_record97_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record114_rec_valid <= main_genericstandalone_rtio_core_sed_record98_rec_valid;
	main_genericstandalone_rtio_core_sed_record114_rec_seqn <= main_genericstandalone_rtio_core_sed_record98_rec_seqn;
	main_genericstandalone_rtio_core_sed_record114_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record98_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record114_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record98_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record114_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record98_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record114_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record98_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record114_rec_payload_address <= main_genericstandalone_rtio_core_sed_record98_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record114_rec_payload_data <= main_genericstandalone_rtio_core_sed_record98_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record115_rec_valid <= main_genericstandalone_rtio_core_sed_record99_rec_valid;
	main_genericstandalone_rtio_core_sed_record115_rec_seqn <= main_genericstandalone_rtio_core_sed_record99_rec_seqn;
	main_genericstandalone_rtio_core_sed_record115_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record99_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record115_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record99_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record115_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record99_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record115_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record99_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record115_rec_payload_address <= main_genericstandalone_rtio_core_sed_record99_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record115_rec_payload_data <= main_genericstandalone_rtio_core_sed_record99_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record124_rec_valid <= main_genericstandalone_rtio_core_sed_record108_rec_valid;
	main_genericstandalone_rtio_core_sed_record124_rec_seqn <= main_genericstandalone_rtio_core_sed_record108_rec_seqn;
	main_genericstandalone_rtio_core_sed_record124_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record108_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record124_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record108_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record124_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record108_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record124_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record108_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record124_rec_payload_address <= main_genericstandalone_rtio_core_sed_record108_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record124_rec_payload_data <= main_genericstandalone_rtio_core_sed_record108_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record125_rec_valid <= main_genericstandalone_rtio_core_sed_record109_rec_valid;
	main_genericstandalone_rtio_core_sed_record125_rec_seqn <= main_genericstandalone_rtio_core_sed_record109_rec_seqn;
	main_genericstandalone_rtio_core_sed_record125_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record109_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record125_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record109_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record125_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record109_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record125_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record109_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record125_rec_payload_address <= main_genericstandalone_rtio_core_sed_record109_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record125_rec_payload_data <= main_genericstandalone_rtio_core_sed_record109_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record126_rec_valid <= main_genericstandalone_rtio_core_sed_record110_rec_valid;
	main_genericstandalone_rtio_core_sed_record126_rec_seqn <= main_genericstandalone_rtio_core_sed_record110_rec_seqn;
	main_genericstandalone_rtio_core_sed_record126_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record110_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record126_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record110_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record126_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record110_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record126_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record110_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record126_rec_payload_address <= main_genericstandalone_rtio_core_sed_record110_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record126_rec_payload_data <= main_genericstandalone_rtio_core_sed_record110_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record127_rec_valid <= main_genericstandalone_rtio_core_sed_record111_rec_valid;
	main_genericstandalone_rtio_core_sed_record127_rec_seqn <= main_genericstandalone_rtio_core_sed_record111_rec_seqn;
	main_genericstandalone_rtio_core_sed_record127_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record111_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record127_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record111_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record127_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record111_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record127_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record111_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record127_rec_payload_address <= main_genericstandalone_rtio_core_sed_record111_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record127_rec_payload_data <= main_genericstandalone_rtio_core_sed_record111_rec_payload_data;
	if (({(~main_genericstandalone_rtio_core_sed_record114_rec_valid), main_genericstandalone_rtio_core_sed_record114_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record116_rec_valid), main_genericstandalone_rtio_core_sed_record116_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record114_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record114_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record116_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record116_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record114_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record116_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record114_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record114_rec_seqn < main_genericstandalone_rtio_core_sed_record116_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record130_rec_valid <= main_genericstandalone_rtio_core_sed_record116_rec_valid;
			main_genericstandalone_rtio_core_sed_record130_rec_seqn <= main_genericstandalone_rtio_core_sed_record116_rec_seqn;
			main_genericstandalone_rtio_core_sed_record130_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record116_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record116_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_address <= main_genericstandalone_rtio_core_sed_record116_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_data <= main_genericstandalone_rtio_core_sed_record116_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record132_rec_valid <= main_genericstandalone_rtio_core_sed_record114_rec_valid;
			main_genericstandalone_rtio_core_sed_record132_rec_seqn <= main_genericstandalone_rtio_core_sed_record114_rec_seqn;
			main_genericstandalone_rtio_core_sed_record132_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record114_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record114_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record114_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record114_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_address <= main_genericstandalone_rtio_core_sed_record114_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_data <= main_genericstandalone_rtio_core_sed_record114_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record130_rec_valid <= main_genericstandalone_rtio_core_sed_record114_rec_valid;
			main_genericstandalone_rtio_core_sed_record130_rec_seqn <= main_genericstandalone_rtio_core_sed_record114_rec_seqn;
			main_genericstandalone_rtio_core_sed_record130_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record114_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record114_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record114_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record114_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_address <= main_genericstandalone_rtio_core_sed_record114_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_data <= main_genericstandalone_rtio_core_sed_record114_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record132_rec_valid <= main_genericstandalone_rtio_core_sed_record116_rec_valid;
			main_genericstandalone_rtio_core_sed_record132_rec_seqn <= main_genericstandalone_rtio_core_sed_record116_rec_seqn;
			main_genericstandalone_rtio_core_sed_record132_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record116_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record116_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_address <= main_genericstandalone_rtio_core_sed_record116_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_data <= main_genericstandalone_rtio_core_sed_record116_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record130_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference50;
		main_genericstandalone_rtio_core_sed_record132_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record114_rec_valid), main_genericstandalone_rtio_core_sed_record114_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record116_rec_valid), main_genericstandalone_rtio_core_sed_record116_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record130_rec_valid <= main_genericstandalone_rtio_core_sed_record114_rec_valid;
			main_genericstandalone_rtio_core_sed_record130_rec_seqn <= main_genericstandalone_rtio_core_sed_record114_rec_seqn;
			main_genericstandalone_rtio_core_sed_record130_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record114_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record114_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record114_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record114_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_address <= main_genericstandalone_rtio_core_sed_record114_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_data <= main_genericstandalone_rtio_core_sed_record114_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record132_rec_valid <= main_genericstandalone_rtio_core_sed_record116_rec_valid;
			main_genericstandalone_rtio_core_sed_record132_rec_seqn <= main_genericstandalone_rtio_core_sed_record116_rec_seqn;
			main_genericstandalone_rtio_core_sed_record132_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record116_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record116_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_address <= main_genericstandalone_rtio_core_sed_record116_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_data <= main_genericstandalone_rtio_core_sed_record116_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record130_rec_valid <= main_genericstandalone_rtio_core_sed_record116_rec_valid;
			main_genericstandalone_rtio_core_sed_record130_rec_seqn <= main_genericstandalone_rtio_core_sed_record116_rec_seqn;
			main_genericstandalone_rtio_core_sed_record130_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record116_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record116_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record116_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record116_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_address <= main_genericstandalone_rtio_core_sed_record116_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record130_rec_payload_data <= main_genericstandalone_rtio_core_sed_record116_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record132_rec_valid <= main_genericstandalone_rtio_core_sed_record114_rec_valid;
			main_genericstandalone_rtio_core_sed_record132_rec_seqn <= main_genericstandalone_rtio_core_sed_record114_rec_seqn;
			main_genericstandalone_rtio_core_sed_record132_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record114_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record114_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record114_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record114_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_address <= main_genericstandalone_rtio_core_sed_record114_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record132_rec_payload_data <= main_genericstandalone_rtio_core_sed_record114_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record115_rec_valid), main_genericstandalone_rtio_core_sed_record115_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record117_rec_valid), main_genericstandalone_rtio_core_sed_record117_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record115_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record115_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record117_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record117_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record115_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record117_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record115_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record115_rec_seqn < main_genericstandalone_rtio_core_sed_record117_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record131_rec_valid <= main_genericstandalone_rtio_core_sed_record117_rec_valid;
			main_genericstandalone_rtio_core_sed_record131_rec_seqn <= main_genericstandalone_rtio_core_sed_record117_rec_seqn;
			main_genericstandalone_rtio_core_sed_record131_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record117_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record117_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_address <= main_genericstandalone_rtio_core_sed_record117_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_data <= main_genericstandalone_rtio_core_sed_record117_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record133_rec_valid <= main_genericstandalone_rtio_core_sed_record115_rec_valid;
			main_genericstandalone_rtio_core_sed_record133_rec_seqn <= main_genericstandalone_rtio_core_sed_record115_rec_seqn;
			main_genericstandalone_rtio_core_sed_record133_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record115_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record115_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record115_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record115_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_address <= main_genericstandalone_rtio_core_sed_record115_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_data <= main_genericstandalone_rtio_core_sed_record115_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record131_rec_valid <= main_genericstandalone_rtio_core_sed_record115_rec_valid;
			main_genericstandalone_rtio_core_sed_record131_rec_seqn <= main_genericstandalone_rtio_core_sed_record115_rec_seqn;
			main_genericstandalone_rtio_core_sed_record131_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record115_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record115_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record115_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record115_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_address <= main_genericstandalone_rtio_core_sed_record115_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_data <= main_genericstandalone_rtio_core_sed_record115_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record133_rec_valid <= main_genericstandalone_rtio_core_sed_record117_rec_valid;
			main_genericstandalone_rtio_core_sed_record133_rec_seqn <= main_genericstandalone_rtio_core_sed_record117_rec_seqn;
			main_genericstandalone_rtio_core_sed_record133_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record117_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record117_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_address <= main_genericstandalone_rtio_core_sed_record117_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_data <= main_genericstandalone_rtio_core_sed_record117_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record131_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference51;
		main_genericstandalone_rtio_core_sed_record133_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record115_rec_valid), main_genericstandalone_rtio_core_sed_record115_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record117_rec_valid), main_genericstandalone_rtio_core_sed_record117_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record131_rec_valid <= main_genericstandalone_rtio_core_sed_record115_rec_valid;
			main_genericstandalone_rtio_core_sed_record131_rec_seqn <= main_genericstandalone_rtio_core_sed_record115_rec_seqn;
			main_genericstandalone_rtio_core_sed_record131_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record115_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record115_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record115_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record115_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_address <= main_genericstandalone_rtio_core_sed_record115_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_data <= main_genericstandalone_rtio_core_sed_record115_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record133_rec_valid <= main_genericstandalone_rtio_core_sed_record117_rec_valid;
			main_genericstandalone_rtio_core_sed_record133_rec_seqn <= main_genericstandalone_rtio_core_sed_record117_rec_seqn;
			main_genericstandalone_rtio_core_sed_record133_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record117_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record117_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_address <= main_genericstandalone_rtio_core_sed_record117_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_data <= main_genericstandalone_rtio_core_sed_record117_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record131_rec_valid <= main_genericstandalone_rtio_core_sed_record117_rec_valid;
			main_genericstandalone_rtio_core_sed_record131_rec_seqn <= main_genericstandalone_rtio_core_sed_record117_rec_seqn;
			main_genericstandalone_rtio_core_sed_record131_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record117_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record117_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record117_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record117_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_address <= main_genericstandalone_rtio_core_sed_record117_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record131_rec_payload_data <= main_genericstandalone_rtio_core_sed_record117_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record133_rec_valid <= main_genericstandalone_rtio_core_sed_record115_rec_valid;
			main_genericstandalone_rtio_core_sed_record133_rec_seqn <= main_genericstandalone_rtio_core_sed_record115_rec_seqn;
			main_genericstandalone_rtio_core_sed_record133_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record115_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record115_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record115_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record115_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_address <= main_genericstandalone_rtio_core_sed_record115_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record133_rec_payload_data <= main_genericstandalone_rtio_core_sed_record115_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record118_rec_valid), main_genericstandalone_rtio_core_sed_record118_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record120_rec_valid), main_genericstandalone_rtio_core_sed_record120_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record118_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record118_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record120_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record120_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record118_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record120_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record118_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record118_rec_seqn < main_genericstandalone_rtio_core_sed_record120_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record134_rec_valid <= main_genericstandalone_rtio_core_sed_record120_rec_valid;
			main_genericstandalone_rtio_core_sed_record134_rec_seqn <= main_genericstandalone_rtio_core_sed_record120_rec_seqn;
			main_genericstandalone_rtio_core_sed_record134_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record120_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record120_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_address <= main_genericstandalone_rtio_core_sed_record120_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_data <= main_genericstandalone_rtio_core_sed_record120_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record136_rec_valid <= main_genericstandalone_rtio_core_sed_record118_rec_valid;
			main_genericstandalone_rtio_core_sed_record136_rec_seqn <= main_genericstandalone_rtio_core_sed_record118_rec_seqn;
			main_genericstandalone_rtio_core_sed_record136_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record118_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record118_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_address <= main_genericstandalone_rtio_core_sed_record118_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_data <= main_genericstandalone_rtio_core_sed_record118_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record134_rec_valid <= main_genericstandalone_rtio_core_sed_record118_rec_valid;
			main_genericstandalone_rtio_core_sed_record134_rec_seqn <= main_genericstandalone_rtio_core_sed_record118_rec_seqn;
			main_genericstandalone_rtio_core_sed_record134_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record118_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record118_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_address <= main_genericstandalone_rtio_core_sed_record118_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_data <= main_genericstandalone_rtio_core_sed_record118_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record136_rec_valid <= main_genericstandalone_rtio_core_sed_record120_rec_valid;
			main_genericstandalone_rtio_core_sed_record136_rec_seqn <= main_genericstandalone_rtio_core_sed_record120_rec_seqn;
			main_genericstandalone_rtio_core_sed_record136_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record120_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record120_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_address <= main_genericstandalone_rtio_core_sed_record120_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_data <= main_genericstandalone_rtio_core_sed_record120_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record134_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference52;
		main_genericstandalone_rtio_core_sed_record136_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record118_rec_valid), main_genericstandalone_rtio_core_sed_record118_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record120_rec_valid), main_genericstandalone_rtio_core_sed_record120_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record134_rec_valid <= main_genericstandalone_rtio_core_sed_record118_rec_valid;
			main_genericstandalone_rtio_core_sed_record134_rec_seqn <= main_genericstandalone_rtio_core_sed_record118_rec_seqn;
			main_genericstandalone_rtio_core_sed_record134_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record118_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record118_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_address <= main_genericstandalone_rtio_core_sed_record118_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_data <= main_genericstandalone_rtio_core_sed_record118_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record136_rec_valid <= main_genericstandalone_rtio_core_sed_record120_rec_valid;
			main_genericstandalone_rtio_core_sed_record136_rec_seqn <= main_genericstandalone_rtio_core_sed_record120_rec_seqn;
			main_genericstandalone_rtio_core_sed_record136_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record120_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record120_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_address <= main_genericstandalone_rtio_core_sed_record120_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_data <= main_genericstandalone_rtio_core_sed_record120_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record134_rec_valid <= main_genericstandalone_rtio_core_sed_record120_rec_valid;
			main_genericstandalone_rtio_core_sed_record134_rec_seqn <= main_genericstandalone_rtio_core_sed_record120_rec_seqn;
			main_genericstandalone_rtio_core_sed_record134_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record120_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record120_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record120_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record120_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_address <= main_genericstandalone_rtio_core_sed_record120_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record134_rec_payload_data <= main_genericstandalone_rtio_core_sed_record120_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record136_rec_valid <= main_genericstandalone_rtio_core_sed_record118_rec_valid;
			main_genericstandalone_rtio_core_sed_record136_rec_seqn <= main_genericstandalone_rtio_core_sed_record118_rec_seqn;
			main_genericstandalone_rtio_core_sed_record136_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record118_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record118_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record118_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record118_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_address <= main_genericstandalone_rtio_core_sed_record118_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record136_rec_payload_data <= main_genericstandalone_rtio_core_sed_record118_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record119_rec_valid), main_genericstandalone_rtio_core_sed_record119_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record121_rec_valid), main_genericstandalone_rtio_core_sed_record121_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record119_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record119_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record121_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record121_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record119_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record121_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record119_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record119_rec_seqn < main_genericstandalone_rtio_core_sed_record121_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record135_rec_valid <= main_genericstandalone_rtio_core_sed_record121_rec_valid;
			main_genericstandalone_rtio_core_sed_record135_rec_seqn <= main_genericstandalone_rtio_core_sed_record121_rec_seqn;
			main_genericstandalone_rtio_core_sed_record135_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record121_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record121_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_address <= main_genericstandalone_rtio_core_sed_record121_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_data <= main_genericstandalone_rtio_core_sed_record121_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record137_rec_valid <= main_genericstandalone_rtio_core_sed_record119_rec_valid;
			main_genericstandalone_rtio_core_sed_record137_rec_seqn <= main_genericstandalone_rtio_core_sed_record119_rec_seqn;
			main_genericstandalone_rtio_core_sed_record137_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record119_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record119_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_address <= main_genericstandalone_rtio_core_sed_record119_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_data <= main_genericstandalone_rtio_core_sed_record119_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record135_rec_valid <= main_genericstandalone_rtio_core_sed_record119_rec_valid;
			main_genericstandalone_rtio_core_sed_record135_rec_seqn <= main_genericstandalone_rtio_core_sed_record119_rec_seqn;
			main_genericstandalone_rtio_core_sed_record135_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record119_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record119_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_address <= main_genericstandalone_rtio_core_sed_record119_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_data <= main_genericstandalone_rtio_core_sed_record119_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record137_rec_valid <= main_genericstandalone_rtio_core_sed_record121_rec_valid;
			main_genericstandalone_rtio_core_sed_record137_rec_seqn <= main_genericstandalone_rtio_core_sed_record121_rec_seqn;
			main_genericstandalone_rtio_core_sed_record137_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record121_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record121_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_address <= main_genericstandalone_rtio_core_sed_record121_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_data <= main_genericstandalone_rtio_core_sed_record121_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record135_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference53;
		main_genericstandalone_rtio_core_sed_record137_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record119_rec_valid), main_genericstandalone_rtio_core_sed_record119_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record121_rec_valid), main_genericstandalone_rtio_core_sed_record121_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record135_rec_valid <= main_genericstandalone_rtio_core_sed_record119_rec_valid;
			main_genericstandalone_rtio_core_sed_record135_rec_seqn <= main_genericstandalone_rtio_core_sed_record119_rec_seqn;
			main_genericstandalone_rtio_core_sed_record135_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record119_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record119_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_address <= main_genericstandalone_rtio_core_sed_record119_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_data <= main_genericstandalone_rtio_core_sed_record119_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record137_rec_valid <= main_genericstandalone_rtio_core_sed_record121_rec_valid;
			main_genericstandalone_rtio_core_sed_record137_rec_seqn <= main_genericstandalone_rtio_core_sed_record121_rec_seqn;
			main_genericstandalone_rtio_core_sed_record137_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record121_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record121_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_address <= main_genericstandalone_rtio_core_sed_record121_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_data <= main_genericstandalone_rtio_core_sed_record121_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record135_rec_valid <= main_genericstandalone_rtio_core_sed_record121_rec_valid;
			main_genericstandalone_rtio_core_sed_record135_rec_seqn <= main_genericstandalone_rtio_core_sed_record121_rec_seqn;
			main_genericstandalone_rtio_core_sed_record135_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record121_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record121_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record121_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record121_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_address <= main_genericstandalone_rtio_core_sed_record121_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record135_rec_payload_data <= main_genericstandalone_rtio_core_sed_record121_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record137_rec_valid <= main_genericstandalone_rtio_core_sed_record119_rec_valid;
			main_genericstandalone_rtio_core_sed_record137_rec_seqn <= main_genericstandalone_rtio_core_sed_record119_rec_seqn;
			main_genericstandalone_rtio_core_sed_record137_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record119_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record119_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record119_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record119_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_address <= main_genericstandalone_rtio_core_sed_record119_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record137_rec_payload_data <= main_genericstandalone_rtio_core_sed_record119_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record122_rec_valid), main_genericstandalone_rtio_core_sed_record122_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record124_rec_valid), main_genericstandalone_rtio_core_sed_record124_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record122_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record122_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record124_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record124_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record122_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record124_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record122_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record122_rec_seqn < main_genericstandalone_rtio_core_sed_record124_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record138_rec_valid <= main_genericstandalone_rtio_core_sed_record124_rec_valid;
			main_genericstandalone_rtio_core_sed_record138_rec_seqn <= main_genericstandalone_rtio_core_sed_record124_rec_seqn;
			main_genericstandalone_rtio_core_sed_record138_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record124_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record124_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record124_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record124_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_address <= main_genericstandalone_rtio_core_sed_record124_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_data <= main_genericstandalone_rtio_core_sed_record124_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record140_rec_valid <= main_genericstandalone_rtio_core_sed_record122_rec_valid;
			main_genericstandalone_rtio_core_sed_record140_rec_seqn <= main_genericstandalone_rtio_core_sed_record122_rec_seqn;
			main_genericstandalone_rtio_core_sed_record140_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record122_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record122_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_address <= main_genericstandalone_rtio_core_sed_record122_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_data <= main_genericstandalone_rtio_core_sed_record122_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record138_rec_valid <= main_genericstandalone_rtio_core_sed_record122_rec_valid;
			main_genericstandalone_rtio_core_sed_record138_rec_seqn <= main_genericstandalone_rtio_core_sed_record122_rec_seqn;
			main_genericstandalone_rtio_core_sed_record138_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record122_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record122_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_address <= main_genericstandalone_rtio_core_sed_record122_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_data <= main_genericstandalone_rtio_core_sed_record122_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record140_rec_valid <= main_genericstandalone_rtio_core_sed_record124_rec_valid;
			main_genericstandalone_rtio_core_sed_record140_rec_seqn <= main_genericstandalone_rtio_core_sed_record124_rec_seqn;
			main_genericstandalone_rtio_core_sed_record140_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record124_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record124_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record124_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record124_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_address <= main_genericstandalone_rtio_core_sed_record124_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_data <= main_genericstandalone_rtio_core_sed_record124_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record138_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference54;
		main_genericstandalone_rtio_core_sed_record140_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record122_rec_valid), main_genericstandalone_rtio_core_sed_record122_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record124_rec_valid), main_genericstandalone_rtio_core_sed_record124_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record138_rec_valid <= main_genericstandalone_rtio_core_sed_record122_rec_valid;
			main_genericstandalone_rtio_core_sed_record138_rec_seqn <= main_genericstandalone_rtio_core_sed_record122_rec_seqn;
			main_genericstandalone_rtio_core_sed_record138_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record122_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record122_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_address <= main_genericstandalone_rtio_core_sed_record122_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_data <= main_genericstandalone_rtio_core_sed_record122_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record140_rec_valid <= main_genericstandalone_rtio_core_sed_record124_rec_valid;
			main_genericstandalone_rtio_core_sed_record140_rec_seqn <= main_genericstandalone_rtio_core_sed_record124_rec_seqn;
			main_genericstandalone_rtio_core_sed_record140_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record124_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record124_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record124_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record124_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_address <= main_genericstandalone_rtio_core_sed_record124_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_data <= main_genericstandalone_rtio_core_sed_record124_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record138_rec_valid <= main_genericstandalone_rtio_core_sed_record124_rec_valid;
			main_genericstandalone_rtio_core_sed_record138_rec_seqn <= main_genericstandalone_rtio_core_sed_record124_rec_seqn;
			main_genericstandalone_rtio_core_sed_record138_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record124_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record124_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record124_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record124_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_address <= main_genericstandalone_rtio_core_sed_record124_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record138_rec_payload_data <= main_genericstandalone_rtio_core_sed_record124_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record140_rec_valid <= main_genericstandalone_rtio_core_sed_record122_rec_valid;
			main_genericstandalone_rtio_core_sed_record140_rec_seqn <= main_genericstandalone_rtio_core_sed_record122_rec_seqn;
			main_genericstandalone_rtio_core_sed_record140_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record122_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record122_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record122_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record122_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_address <= main_genericstandalone_rtio_core_sed_record122_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record140_rec_payload_data <= main_genericstandalone_rtio_core_sed_record122_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record123_rec_valid), main_genericstandalone_rtio_core_sed_record123_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record125_rec_valid), main_genericstandalone_rtio_core_sed_record125_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record123_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record123_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record125_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record125_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record123_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record125_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record123_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record123_rec_seqn < main_genericstandalone_rtio_core_sed_record125_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record139_rec_valid <= main_genericstandalone_rtio_core_sed_record125_rec_valid;
			main_genericstandalone_rtio_core_sed_record139_rec_seqn <= main_genericstandalone_rtio_core_sed_record125_rec_seqn;
			main_genericstandalone_rtio_core_sed_record139_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record125_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record125_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record125_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record125_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_address <= main_genericstandalone_rtio_core_sed_record125_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_data <= main_genericstandalone_rtio_core_sed_record125_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record141_rec_valid <= main_genericstandalone_rtio_core_sed_record123_rec_valid;
			main_genericstandalone_rtio_core_sed_record141_rec_seqn <= main_genericstandalone_rtio_core_sed_record123_rec_seqn;
			main_genericstandalone_rtio_core_sed_record141_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record123_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record123_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_address <= main_genericstandalone_rtio_core_sed_record123_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_data <= main_genericstandalone_rtio_core_sed_record123_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record139_rec_valid <= main_genericstandalone_rtio_core_sed_record123_rec_valid;
			main_genericstandalone_rtio_core_sed_record139_rec_seqn <= main_genericstandalone_rtio_core_sed_record123_rec_seqn;
			main_genericstandalone_rtio_core_sed_record139_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record123_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record123_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_address <= main_genericstandalone_rtio_core_sed_record123_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_data <= main_genericstandalone_rtio_core_sed_record123_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record141_rec_valid <= main_genericstandalone_rtio_core_sed_record125_rec_valid;
			main_genericstandalone_rtio_core_sed_record141_rec_seqn <= main_genericstandalone_rtio_core_sed_record125_rec_seqn;
			main_genericstandalone_rtio_core_sed_record141_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record125_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record125_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record125_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record125_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_address <= main_genericstandalone_rtio_core_sed_record125_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_data <= main_genericstandalone_rtio_core_sed_record125_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record139_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference55;
		main_genericstandalone_rtio_core_sed_record141_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record123_rec_valid), main_genericstandalone_rtio_core_sed_record123_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record125_rec_valid), main_genericstandalone_rtio_core_sed_record125_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record139_rec_valid <= main_genericstandalone_rtio_core_sed_record123_rec_valid;
			main_genericstandalone_rtio_core_sed_record139_rec_seqn <= main_genericstandalone_rtio_core_sed_record123_rec_seqn;
			main_genericstandalone_rtio_core_sed_record139_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record123_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record123_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_address <= main_genericstandalone_rtio_core_sed_record123_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_data <= main_genericstandalone_rtio_core_sed_record123_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record141_rec_valid <= main_genericstandalone_rtio_core_sed_record125_rec_valid;
			main_genericstandalone_rtio_core_sed_record141_rec_seqn <= main_genericstandalone_rtio_core_sed_record125_rec_seqn;
			main_genericstandalone_rtio_core_sed_record141_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record125_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record125_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record125_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record125_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_address <= main_genericstandalone_rtio_core_sed_record125_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_data <= main_genericstandalone_rtio_core_sed_record125_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record139_rec_valid <= main_genericstandalone_rtio_core_sed_record125_rec_valid;
			main_genericstandalone_rtio_core_sed_record139_rec_seqn <= main_genericstandalone_rtio_core_sed_record125_rec_seqn;
			main_genericstandalone_rtio_core_sed_record139_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record125_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record125_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record125_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record125_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_address <= main_genericstandalone_rtio_core_sed_record125_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record139_rec_payload_data <= main_genericstandalone_rtio_core_sed_record125_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record141_rec_valid <= main_genericstandalone_rtio_core_sed_record123_rec_valid;
			main_genericstandalone_rtio_core_sed_record141_rec_seqn <= main_genericstandalone_rtio_core_sed_record123_rec_seqn;
			main_genericstandalone_rtio_core_sed_record141_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record123_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record123_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record123_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record123_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_address <= main_genericstandalone_rtio_core_sed_record123_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record141_rec_payload_data <= main_genericstandalone_rtio_core_sed_record123_rec_payload_data;
		end
	end
	main_genericstandalone_rtio_core_sed_record128_rec_valid <= main_genericstandalone_rtio_core_sed_record112_rec_valid;
	main_genericstandalone_rtio_core_sed_record128_rec_seqn <= main_genericstandalone_rtio_core_sed_record112_rec_seqn;
	main_genericstandalone_rtio_core_sed_record128_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record112_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record128_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record112_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record128_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record112_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record128_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record112_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record128_rec_payload_address <= main_genericstandalone_rtio_core_sed_record112_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record128_rec_payload_data <= main_genericstandalone_rtio_core_sed_record112_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record129_rec_valid <= main_genericstandalone_rtio_core_sed_record113_rec_valid;
	main_genericstandalone_rtio_core_sed_record129_rec_seqn <= main_genericstandalone_rtio_core_sed_record113_rec_seqn;
	main_genericstandalone_rtio_core_sed_record129_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record113_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record129_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record113_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record129_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record113_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record129_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record113_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record129_rec_payload_address <= main_genericstandalone_rtio_core_sed_record113_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record129_rec_payload_data <= main_genericstandalone_rtio_core_sed_record113_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record142_rec_valid <= main_genericstandalone_rtio_core_sed_record126_rec_valid;
	main_genericstandalone_rtio_core_sed_record142_rec_seqn <= main_genericstandalone_rtio_core_sed_record126_rec_seqn;
	main_genericstandalone_rtio_core_sed_record142_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record126_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record142_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record126_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record142_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record126_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record142_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record126_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record142_rec_payload_address <= main_genericstandalone_rtio_core_sed_record126_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record142_rec_payload_data <= main_genericstandalone_rtio_core_sed_record126_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record143_rec_valid <= main_genericstandalone_rtio_core_sed_record127_rec_valid;
	main_genericstandalone_rtio_core_sed_record143_rec_seqn <= main_genericstandalone_rtio_core_sed_record127_rec_seqn;
	main_genericstandalone_rtio_core_sed_record143_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record127_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record143_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record127_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record143_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record127_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record143_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record127_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record143_rec_payload_address <= main_genericstandalone_rtio_core_sed_record127_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record143_rec_payload_data <= main_genericstandalone_rtio_core_sed_record127_rec_payload_data;
	if (({(~main_genericstandalone_rtio_core_sed_record129_rec_valid), main_genericstandalone_rtio_core_sed_record129_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record130_rec_valid), main_genericstandalone_rtio_core_sed_record130_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record129_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record129_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record130_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record130_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record129_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record130_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record129_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record129_rec_seqn < main_genericstandalone_rtio_core_sed_record130_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record145_rec_valid <= main_genericstandalone_rtio_core_sed_record130_rec_valid;
			main_genericstandalone_rtio_core_sed_record145_rec_seqn <= main_genericstandalone_rtio_core_sed_record130_rec_seqn;
			main_genericstandalone_rtio_core_sed_record145_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record130_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record145_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record130_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_address <= main_genericstandalone_rtio_core_sed_record130_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_data <= main_genericstandalone_rtio_core_sed_record130_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record146_rec_valid <= main_genericstandalone_rtio_core_sed_record129_rec_valid;
			main_genericstandalone_rtio_core_sed_record146_rec_seqn <= main_genericstandalone_rtio_core_sed_record129_rec_seqn;
			main_genericstandalone_rtio_core_sed_record146_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record129_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record146_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record129_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record129_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record129_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_address <= main_genericstandalone_rtio_core_sed_record129_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_data <= main_genericstandalone_rtio_core_sed_record129_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record145_rec_valid <= main_genericstandalone_rtio_core_sed_record129_rec_valid;
			main_genericstandalone_rtio_core_sed_record145_rec_seqn <= main_genericstandalone_rtio_core_sed_record129_rec_seqn;
			main_genericstandalone_rtio_core_sed_record145_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record129_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record145_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record129_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record129_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record129_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_address <= main_genericstandalone_rtio_core_sed_record129_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_data <= main_genericstandalone_rtio_core_sed_record129_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record146_rec_valid <= main_genericstandalone_rtio_core_sed_record130_rec_valid;
			main_genericstandalone_rtio_core_sed_record146_rec_seqn <= main_genericstandalone_rtio_core_sed_record130_rec_seqn;
			main_genericstandalone_rtio_core_sed_record146_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record130_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record146_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record130_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_address <= main_genericstandalone_rtio_core_sed_record130_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_data <= main_genericstandalone_rtio_core_sed_record130_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record145_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record145_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference56;
		main_genericstandalone_rtio_core_sed_record146_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record129_rec_valid), main_genericstandalone_rtio_core_sed_record129_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record130_rec_valid), main_genericstandalone_rtio_core_sed_record130_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record145_rec_valid <= main_genericstandalone_rtio_core_sed_record129_rec_valid;
			main_genericstandalone_rtio_core_sed_record145_rec_seqn <= main_genericstandalone_rtio_core_sed_record129_rec_seqn;
			main_genericstandalone_rtio_core_sed_record145_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record129_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record145_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record129_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record129_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record129_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_address <= main_genericstandalone_rtio_core_sed_record129_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_data <= main_genericstandalone_rtio_core_sed_record129_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record146_rec_valid <= main_genericstandalone_rtio_core_sed_record130_rec_valid;
			main_genericstandalone_rtio_core_sed_record146_rec_seqn <= main_genericstandalone_rtio_core_sed_record130_rec_seqn;
			main_genericstandalone_rtio_core_sed_record146_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record130_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record146_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record130_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_address <= main_genericstandalone_rtio_core_sed_record130_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_data <= main_genericstandalone_rtio_core_sed_record130_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record145_rec_valid <= main_genericstandalone_rtio_core_sed_record130_rec_valid;
			main_genericstandalone_rtio_core_sed_record145_rec_seqn <= main_genericstandalone_rtio_core_sed_record130_rec_seqn;
			main_genericstandalone_rtio_core_sed_record145_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record130_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record145_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record130_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record130_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record130_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_address <= main_genericstandalone_rtio_core_sed_record130_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record145_rec_payload_data <= main_genericstandalone_rtio_core_sed_record130_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record146_rec_valid <= main_genericstandalone_rtio_core_sed_record129_rec_valid;
			main_genericstandalone_rtio_core_sed_record146_rec_seqn <= main_genericstandalone_rtio_core_sed_record129_rec_seqn;
			main_genericstandalone_rtio_core_sed_record146_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record129_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record146_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record129_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record129_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record129_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_address <= main_genericstandalone_rtio_core_sed_record129_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record146_rec_payload_data <= main_genericstandalone_rtio_core_sed_record129_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record131_rec_valid), main_genericstandalone_rtio_core_sed_record131_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record132_rec_valid), main_genericstandalone_rtio_core_sed_record132_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record131_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record131_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record132_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record132_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record131_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record132_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record131_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record131_rec_seqn < main_genericstandalone_rtio_core_sed_record132_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record147_rec_valid <= main_genericstandalone_rtio_core_sed_record132_rec_valid;
			main_genericstandalone_rtio_core_sed_record147_rec_seqn <= main_genericstandalone_rtio_core_sed_record132_rec_seqn;
			main_genericstandalone_rtio_core_sed_record147_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record132_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record147_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record132_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_address <= main_genericstandalone_rtio_core_sed_record132_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_data <= main_genericstandalone_rtio_core_sed_record132_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record148_rec_valid <= main_genericstandalone_rtio_core_sed_record131_rec_valid;
			main_genericstandalone_rtio_core_sed_record148_rec_seqn <= main_genericstandalone_rtio_core_sed_record131_rec_seqn;
			main_genericstandalone_rtio_core_sed_record148_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record131_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record148_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record131_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_address <= main_genericstandalone_rtio_core_sed_record131_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_data <= main_genericstandalone_rtio_core_sed_record131_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record147_rec_valid <= main_genericstandalone_rtio_core_sed_record131_rec_valid;
			main_genericstandalone_rtio_core_sed_record147_rec_seqn <= main_genericstandalone_rtio_core_sed_record131_rec_seqn;
			main_genericstandalone_rtio_core_sed_record147_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record131_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record147_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record131_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_address <= main_genericstandalone_rtio_core_sed_record131_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_data <= main_genericstandalone_rtio_core_sed_record131_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record148_rec_valid <= main_genericstandalone_rtio_core_sed_record132_rec_valid;
			main_genericstandalone_rtio_core_sed_record148_rec_seqn <= main_genericstandalone_rtio_core_sed_record132_rec_seqn;
			main_genericstandalone_rtio_core_sed_record148_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record132_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record148_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record132_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_address <= main_genericstandalone_rtio_core_sed_record132_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_data <= main_genericstandalone_rtio_core_sed_record132_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record147_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record147_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference57;
		main_genericstandalone_rtio_core_sed_record148_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record131_rec_valid), main_genericstandalone_rtio_core_sed_record131_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record132_rec_valid), main_genericstandalone_rtio_core_sed_record132_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record147_rec_valid <= main_genericstandalone_rtio_core_sed_record131_rec_valid;
			main_genericstandalone_rtio_core_sed_record147_rec_seqn <= main_genericstandalone_rtio_core_sed_record131_rec_seqn;
			main_genericstandalone_rtio_core_sed_record147_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record131_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record147_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record131_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_address <= main_genericstandalone_rtio_core_sed_record131_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_data <= main_genericstandalone_rtio_core_sed_record131_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record148_rec_valid <= main_genericstandalone_rtio_core_sed_record132_rec_valid;
			main_genericstandalone_rtio_core_sed_record148_rec_seqn <= main_genericstandalone_rtio_core_sed_record132_rec_seqn;
			main_genericstandalone_rtio_core_sed_record148_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record132_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record148_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record132_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_address <= main_genericstandalone_rtio_core_sed_record132_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_data <= main_genericstandalone_rtio_core_sed_record132_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record147_rec_valid <= main_genericstandalone_rtio_core_sed_record132_rec_valid;
			main_genericstandalone_rtio_core_sed_record147_rec_seqn <= main_genericstandalone_rtio_core_sed_record132_rec_seqn;
			main_genericstandalone_rtio_core_sed_record147_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record132_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record147_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record132_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record132_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record132_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_address <= main_genericstandalone_rtio_core_sed_record132_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record147_rec_payload_data <= main_genericstandalone_rtio_core_sed_record132_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record148_rec_valid <= main_genericstandalone_rtio_core_sed_record131_rec_valid;
			main_genericstandalone_rtio_core_sed_record148_rec_seqn <= main_genericstandalone_rtio_core_sed_record131_rec_seqn;
			main_genericstandalone_rtio_core_sed_record148_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record131_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record148_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record131_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record131_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record131_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_address <= main_genericstandalone_rtio_core_sed_record131_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record148_rec_payload_data <= main_genericstandalone_rtio_core_sed_record131_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record133_rec_valid), main_genericstandalone_rtio_core_sed_record133_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record134_rec_valid), main_genericstandalone_rtio_core_sed_record134_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record133_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record133_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record134_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record134_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record133_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record134_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record133_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record133_rec_seqn < main_genericstandalone_rtio_core_sed_record134_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record149_rec_valid <= main_genericstandalone_rtio_core_sed_record134_rec_valid;
			main_genericstandalone_rtio_core_sed_record149_rec_seqn <= main_genericstandalone_rtio_core_sed_record134_rec_seqn;
			main_genericstandalone_rtio_core_sed_record149_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record134_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record149_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record134_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_address <= main_genericstandalone_rtio_core_sed_record134_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_data <= main_genericstandalone_rtio_core_sed_record134_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record150_rec_valid <= main_genericstandalone_rtio_core_sed_record133_rec_valid;
			main_genericstandalone_rtio_core_sed_record150_rec_seqn <= main_genericstandalone_rtio_core_sed_record133_rec_seqn;
			main_genericstandalone_rtio_core_sed_record150_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record133_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record150_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record133_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_address <= main_genericstandalone_rtio_core_sed_record133_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_data <= main_genericstandalone_rtio_core_sed_record133_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record149_rec_valid <= main_genericstandalone_rtio_core_sed_record133_rec_valid;
			main_genericstandalone_rtio_core_sed_record149_rec_seqn <= main_genericstandalone_rtio_core_sed_record133_rec_seqn;
			main_genericstandalone_rtio_core_sed_record149_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record133_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record149_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record133_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_address <= main_genericstandalone_rtio_core_sed_record133_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_data <= main_genericstandalone_rtio_core_sed_record133_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record150_rec_valid <= main_genericstandalone_rtio_core_sed_record134_rec_valid;
			main_genericstandalone_rtio_core_sed_record150_rec_seqn <= main_genericstandalone_rtio_core_sed_record134_rec_seqn;
			main_genericstandalone_rtio_core_sed_record150_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record134_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record150_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record134_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_address <= main_genericstandalone_rtio_core_sed_record134_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_data <= main_genericstandalone_rtio_core_sed_record134_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record149_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record149_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference58;
		main_genericstandalone_rtio_core_sed_record150_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record133_rec_valid), main_genericstandalone_rtio_core_sed_record133_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record134_rec_valid), main_genericstandalone_rtio_core_sed_record134_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record149_rec_valid <= main_genericstandalone_rtio_core_sed_record133_rec_valid;
			main_genericstandalone_rtio_core_sed_record149_rec_seqn <= main_genericstandalone_rtio_core_sed_record133_rec_seqn;
			main_genericstandalone_rtio_core_sed_record149_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record133_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record149_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record133_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_address <= main_genericstandalone_rtio_core_sed_record133_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_data <= main_genericstandalone_rtio_core_sed_record133_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record150_rec_valid <= main_genericstandalone_rtio_core_sed_record134_rec_valid;
			main_genericstandalone_rtio_core_sed_record150_rec_seqn <= main_genericstandalone_rtio_core_sed_record134_rec_seqn;
			main_genericstandalone_rtio_core_sed_record150_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record134_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record150_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record134_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_address <= main_genericstandalone_rtio_core_sed_record134_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_data <= main_genericstandalone_rtio_core_sed_record134_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record149_rec_valid <= main_genericstandalone_rtio_core_sed_record134_rec_valid;
			main_genericstandalone_rtio_core_sed_record149_rec_seqn <= main_genericstandalone_rtio_core_sed_record134_rec_seqn;
			main_genericstandalone_rtio_core_sed_record149_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record134_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record149_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record134_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record134_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record134_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_address <= main_genericstandalone_rtio_core_sed_record134_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record149_rec_payload_data <= main_genericstandalone_rtio_core_sed_record134_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record150_rec_valid <= main_genericstandalone_rtio_core_sed_record133_rec_valid;
			main_genericstandalone_rtio_core_sed_record150_rec_seqn <= main_genericstandalone_rtio_core_sed_record133_rec_seqn;
			main_genericstandalone_rtio_core_sed_record150_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record133_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record150_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record133_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record133_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record133_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_address <= main_genericstandalone_rtio_core_sed_record133_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record150_rec_payload_data <= main_genericstandalone_rtio_core_sed_record133_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record135_rec_valid), main_genericstandalone_rtio_core_sed_record135_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record136_rec_valid), main_genericstandalone_rtio_core_sed_record136_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record135_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record135_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record136_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record136_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record135_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record136_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record135_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record135_rec_seqn < main_genericstandalone_rtio_core_sed_record136_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record151_rec_valid <= main_genericstandalone_rtio_core_sed_record136_rec_valid;
			main_genericstandalone_rtio_core_sed_record151_rec_seqn <= main_genericstandalone_rtio_core_sed_record136_rec_seqn;
			main_genericstandalone_rtio_core_sed_record151_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record136_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record151_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record136_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_address <= main_genericstandalone_rtio_core_sed_record136_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_data <= main_genericstandalone_rtio_core_sed_record136_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record152_rec_valid <= main_genericstandalone_rtio_core_sed_record135_rec_valid;
			main_genericstandalone_rtio_core_sed_record152_rec_seqn <= main_genericstandalone_rtio_core_sed_record135_rec_seqn;
			main_genericstandalone_rtio_core_sed_record152_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record135_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record152_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record135_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_address <= main_genericstandalone_rtio_core_sed_record135_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_data <= main_genericstandalone_rtio_core_sed_record135_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record151_rec_valid <= main_genericstandalone_rtio_core_sed_record135_rec_valid;
			main_genericstandalone_rtio_core_sed_record151_rec_seqn <= main_genericstandalone_rtio_core_sed_record135_rec_seqn;
			main_genericstandalone_rtio_core_sed_record151_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record135_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record151_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record135_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_address <= main_genericstandalone_rtio_core_sed_record135_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_data <= main_genericstandalone_rtio_core_sed_record135_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record152_rec_valid <= main_genericstandalone_rtio_core_sed_record136_rec_valid;
			main_genericstandalone_rtio_core_sed_record152_rec_seqn <= main_genericstandalone_rtio_core_sed_record136_rec_seqn;
			main_genericstandalone_rtio_core_sed_record152_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record136_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record152_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record136_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_address <= main_genericstandalone_rtio_core_sed_record136_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_data <= main_genericstandalone_rtio_core_sed_record136_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record151_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record151_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference59;
		main_genericstandalone_rtio_core_sed_record152_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record135_rec_valid), main_genericstandalone_rtio_core_sed_record135_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record136_rec_valid), main_genericstandalone_rtio_core_sed_record136_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record151_rec_valid <= main_genericstandalone_rtio_core_sed_record135_rec_valid;
			main_genericstandalone_rtio_core_sed_record151_rec_seqn <= main_genericstandalone_rtio_core_sed_record135_rec_seqn;
			main_genericstandalone_rtio_core_sed_record151_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record135_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record151_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record135_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_address <= main_genericstandalone_rtio_core_sed_record135_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_data <= main_genericstandalone_rtio_core_sed_record135_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record152_rec_valid <= main_genericstandalone_rtio_core_sed_record136_rec_valid;
			main_genericstandalone_rtio_core_sed_record152_rec_seqn <= main_genericstandalone_rtio_core_sed_record136_rec_seqn;
			main_genericstandalone_rtio_core_sed_record152_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record136_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record152_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record136_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_address <= main_genericstandalone_rtio_core_sed_record136_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_data <= main_genericstandalone_rtio_core_sed_record136_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record151_rec_valid <= main_genericstandalone_rtio_core_sed_record136_rec_valid;
			main_genericstandalone_rtio_core_sed_record151_rec_seqn <= main_genericstandalone_rtio_core_sed_record136_rec_seqn;
			main_genericstandalone_rtio_core_sed_record151_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record136_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record151_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record136_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record136_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record136_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_address <= main_genericstandalone_rtio_core_sed_record136_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record151_rec_payload_data <= main_genericstandalone_rtio_core_sed_record136_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record152_rec_valid <= main_genericstandalone_rtio_core_sed_record135_rec_valid;
			main_genericstandalone_rtio_core_sed_record152_rec_seqn <= main_genericstandalone_rtio_core_sed_record135_rec_seqn;
			main_genericstandalone_rtio_core_sed_record152_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record135_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record152_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record135_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record135_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record135_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_address <= main_genericstandalone_rtio_core_sed_record135_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record152_rec_payload_data <= main_genericstandalone_rtio_core_sed_record135_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record137_rec_valid), main_genericstandalone_rtio_core_sed_record137_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record138_rec_valid), main_genericstandalone_rtio_core_sed_record138_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record137_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record137_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record138_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record138_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record137_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record138_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record137_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record137_rec_seqn < main_genericstandalone_rtio_core_sed_record138_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record153_rec_valid <= main_genericstandalone_rtio_core_sed_record138_rec_valid;
			main_genericstandalone_rtio_core_sed_record153_rec_seqn <= main_genericstandalone_rtio_core_sed_record138_rec_seqn;
			main_genericstandalone_rtio_core_sed_record153_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record138_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record153_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record138_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_address <= main_genericstandalone_rtio_core_sed_record138_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_data <= main_genericstandalone_rtio_core_sed_record138_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record154_rec_valid <= main_genericstandalone_rtio_core_sed_record137_rec_valid;
			main_genericstandalone_rtio_core_sed_record154_rec_seqn <= main_genericstandalone_rtio_core_sed_record137_rec_seqn;
			main_genericstandalone_rtio_core_sed_record154_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record137_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record154_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record137_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_address <= main_genericstandalone_rtio_core_sed_record137_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_data <= main_genericstandalone_rtio_core_sed_record137_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record153_rec_valid <= main_genericstandalone_rtio_core_sed_record137_rec_valid;
			main_genericstandalone_rtio_core_sed_record153_rec_seqn <= main_genericstandalone_rtio_core_sed_record137_rec_seqn;
			main_genericstandalone_rtio_core_sed_record153_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record137_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record153_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record137_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_address <= main_genericstandalone_rtio_core_sed_record137_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_data <= main_genericstandalone_rtio_core_sed_record137_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record154_rec_valid <= main_genericstandalone_rtio_core_sed_record138_rec_valid;
			main_genericstandalone_rtio_core_sed_record154_rec_seqn <= main_genericstandalone_rtio_core_sed_record138_rec_seqn;
			main_genericstandalone_rtio_core_sed_record154_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record138_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record154_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record138_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_address <= main_genericstandalone_rtio_core_sed_record138_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_data <= main_genericstandalone_rtio_core_sed_record138_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record153_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record153_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference60;
		main_genericstandalone_rtio_core_sed_record154_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record137_rec_valid), main_genericstandalone_rtio_core_sed_record137_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record138_rec_valid), main_genericstandalone_rtio_core_sed_record138_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record153_rec_valid <= main_genericstandalone_rtio_core_sed_record137_rec_valid;
			main_genericstandalone_rtio_core_sed_record153_rec_seqn <= main_genericstandalone_rtio_core_sed_record137_rec_seqn;
			main_genericstandalone_rtio_core_sed_record153_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record137_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record153_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record137_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_address <= main_genericstandalone_rtio_core_sed_record137_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_data <= main_genericstandalone_rtio_core_sed_record137_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record154_rec_valid <= main_genericstandalone_rtio_core_sed_record138_rec_valid;
			main_genericstandalone_rtio_core_sed_record154_rec_seqn <= main_genericstandalone_rtio_core_sed_record138_rec_seqn;
			main_genericstandalone_rtio_core_sed_record154_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record138_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record154_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record138_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_address <= main_genericstandalone_rtio_core_sed_record138_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_data <= main_genericstandalone_rtio_core_sed_record138_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record153_rec_valid <= main_genericstandalone_rtio_core_sed_record138_rec_valid;
			main_genericstandalone_rtio_core_sed_record153_rec_seqn <= main_genericstandalone_rtio_core_sed_record138_rec_seqn;
			main_genericstandalone_rtio_core_sed_record153_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record138_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record153_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record138_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record138_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record138_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_address <= main_genericstandalone_rtio_core_sed_record138_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record153_rec_payload_data <= main_genericstandalone_rtio_core_sed_record138_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record154_rec_valid <= main_genericstandalone_rtio_core_sed_record137_rec_valid;
			main_genericstandalone_rtio_core_sed_record154_rec_seqn <= main_genericstandalone_rtio_core_sed_record137_rec_seqn;
			main_genericstandalone_rtio_core_sed_record154_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record137_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record154_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record137_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record137_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record137_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_address <= main_genericstandalone_rtio_core_sed_record137_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record154_rec_payload_data <= main_genericstandalone_rtio_core_sed_record137_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record139_rec_valid), main_genericstandalone_rtio_core_sed_record139_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record140_rec_valid), main_genericstandalone_rtio_core_sed_record140_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record139_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record139_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record140_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record140_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record139_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record140_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record139_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record139_rec_seqn < main_genericstandalone_rtio_core_sed_record140_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record155_rec_valid <= main_genericstandalone_rtio_core_sed_record140_rec_valid;
			main_genericstandalone_rtio_core_sed_record155_rec_seqn <= main_genericstandalone_rtio_core_sed_record140_rec_seqn;
			main_genericstandalone_rtio_core_sed_record155_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record140_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record155_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record140_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_address <= main_genericstandalone_rtio_core_sed_record140_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_data <= main_genericstandalone_rtio_core_sed_record140_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record156_rec_valid <= main_genericstandalone_rtio_core_sed_record139_rec_valid;
			main_genericstandalone_rtio_core_sed_record156_rec_seqn <= main_genericstandalone_rtio_core_sed_record139_rec_seqn;
			main_genericstandalone_rtio_core_sed_record156_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record139_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record156_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record139_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_address <= main_genericstandalone_rtio_core_sed_record139_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_data <= main_genericstandalone_rtio_core_sed_record139_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record155_rec_valid <= main_genericstandalone_rtio_core_sed_record139_rec_valid;
			main_genericstandalone_rtio_core_sed_record155_rec_seqn <= main_genericstandalone_rtio_core_sed_record139_rec_seqn;
			main_genericstandalone_rtio_core_sed_record155_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record139_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record155_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record139_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_address <= main_genericstandalone_rtio_core_sed_record139_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_data <= main_genericstandalone_rtio_core_sed_record139_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record156_rec_valid <= main_genericstandalone_rtio_core_sed_record140_rec_valid;
			main_genericstandalone_rtio_core_sed_record156_rec_seqn <= main_genericstandalone_rtio_core_sed_record140_rec_seqn;
			main_genericstandalone_rtio_core_sed_record156_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record140_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record156_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record140_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_address <= main_genericstandalone_rtio_core_sed_record140_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_data <= main_genericstandalone_rtio_core_sed_record140_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record155_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record155_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference61;
		main_genericstandalone_rtio_core_sed_record156_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record139_rec_valid), main_genericstandalone_rtio_core_sed_record139_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record140_rec_valid), main_genericstandalone_rtio_core_sed_record140_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record155_rec_valid <= main_genericstandalone_rtio_core_sed_record139_rec_valid;
			main_genericstandalone_rtio_core_sed_record155_rec_seqn <= main_genericstandalone_rtio_core_sed_record139_rec_seqn;
			main_genericstandalone_rtio_core_sed_record155_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record139_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record155_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record139_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_address <= main_genericstandalone_rtio_core_sed_record139_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_data <= main_genericstandalone_rtio_core_sed_record139_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record156_rec_valid <= main_genericstandalone_rtio_core_sed_record140_rec_valid;
			main_genericstandalone_rtio_core_sed_record156_rec_seqn <= main_genericstandalone_rtio_core_sed_record140_rec_seqn;
			main_genericstandalone_rtio_core_sed_record156_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record140_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record156_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record140_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_address <= main_genericstandalone_rtio_core_sed_record140_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_data <= main_genericstandalone_rtio_core_sed_record140_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record155_rec_valid <= main_genericstandalone_rtio_core_sed_record140_rec_valid;
			main_genericstandalone_rtio_core_sed_record155_rec_seqn <= main_genericstandalone_rtio_core_sed_record140_rec_seqn;
			main_genericstandalone_rtio_core_sed_record155_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record140_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record155_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record140_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record140_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record140_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_address <= main_genericstandalone_rtio_core_sed_record140_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record155_rec_payload_data <= main_genericstandalone_rtio_core_sed_record140_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record156_rec_valid <= main_genericstandalone_rtio_core_sed_record139_rec_valid;
			main_genericstandalone_rtio_core_sed_record156_rec_seqn <= main_genericstandalone_rtio_core_sed_record139_rec_seqn;
			main_genericstandalone_rtio_core_sed_record156_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record139_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record156_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record139_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record139_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record139_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_address <= main_genericstandalone_rtio_core_sed_record139_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record156_rec_payload_data <= main_genericstandalone_rtio_core_sed_record139_rec_payload_data;
		end
	end
	if (({(~main_genericstandalone_rtio_core_sed_record141_rec_valid), main_genericstandalone_rtio_core_sed_record141_rec_payload_channel} == {(~main_genericstandalone_rtio_core_sed_record142_rec_valid), main_genericstandalone_rtio_core_sed_record142_rec_payload_channel})) begin
		if (((((main_genericstandalone_rtio_core_sed_record141_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record141_rec_seqn[12]) & (main_genericstandalone_rtio_core_sed_record142_rec_seqn[11] == main_genericstandalone_rtio_core_sed_record142_rec_seqn[12])) & (main_genericstandalone_rtio_core_sed_record141_rec_seqn[12] != main_genericstandalone_rtio_core_sed_record142_rec_seqn[12])) ? main_genericstandalone_rtio_core_sed_record141_rec_seqn[12] : (main_genericstandalone_rtio_core_sed_record141_rec_seqn < main_genericstandalone_rtio_core_sed_record142_rec_seqn))) begin
			main_genericstandalone_rtio_core_sed_record157_rec_valid <= main_genericstandalone_rtio_core_sed_record142_rec_valid;
			main_genericstandalone_rtio_core_sed_record157_rec_seqn <= main_genericstandalone_rtio_core_sed_record142_rec_seqn;
			main_genericstandalone_rtio_core_sed_record157_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record142_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record157_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record142_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record142_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record142_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_address <= main_genericstandalone_rtio_core_sed_record142_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_data <= main_genericstandalone_rtio_core_sed_record142_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record158_rec_valid <= main_genericstandalone_rtio_core_sed_record141_rec_valid;
			main_genericstandalone_rtio_core_sed_record158_rec_seqn <= main_genericstandalone_rtio_core_sed_record141_rec_seqn;
			main_genericstandalone_rtio_core_sed_record158_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record141_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record158_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record141_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_address <= main_genericstandalone_rtio_core_sed_record141_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_data <= main_genericstandalone_rtio_core_sed_record141_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record157_rec_valid <= main_genericstandalone_rtio_core_sed_record141_rec_valid;
			main_genericstandalone_rtio_core_sed_record157_rec_seqn <= main_genericstandalone_rtio_core_sed_record141_rec_seqn;
			main_genericstandalone_rtio_core_sed_record157_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record141_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record157_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record141_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_address <= main_genericstandalone_rtio_core_sed_record141_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_data <= main_genericstandalone_rtio_core_sed_record141_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record158_rec_valid <= main_genericstandalone_rtio_core_sed_record142_rec_valid;
			main_genericstandalone_rtio_core_sed_record158_rec_seqn <= main_genericstandalone_rtio_core_sed_record142_rec_seqn;
			main_genericstandalone_rtio_core_sed_record158_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record142_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record158_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record142_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record142_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record142_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_address <= main_genericstandalone_rtio_core_sed_record142_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_data <= main_genericstandalone_rtio_core_sed_record142_rec_payload_data;
		end
		main_genericstandalone_rtio_core_sed_record157_rec_replace_occured <= 1'd1;
		main_genericstandalone_rtio_core_sed_record157_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_nondata_difference62;
		main_genericstandalone_rtio_core_sed_record158_rec_valid <= 1'd0;
	end else begin
		if (({(~main_genericstandalone_rtio_core_sed_record141_rec_valid), main_genericstandalone_rtio_core_sed_record141_rec_payload_channel} < {(~main_genericstandalone_rtio_core_sed_record142_rec_valid), main_genericstandalone_rtio_core_sed_record142_rec_payload_channel})) begin
			main_genericstandalone_rtio_core_sed_record157_rec_valid <= main_genericstandalone_rtio_core_sed_record141_rec_valid;
			main_genericstandalone_rtio_core_sed_record157_rec_seqn <= main_genericstandalone_rtio_core_sed_record141_rec_seqn;
			main_genericstandalone_rtio_core_sed_record157_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record141_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record157_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record141_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_address <= main_genericstandalone_rtio_core_sed_record141_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_data <= main_genericstandalone_rtio_core_sed_record141_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record158_rec_valid <= main_genericstandalone_rtio_core_sed_record142_rec_valid;
			main_genericstandalone_rtio_core_sed_record158_rec_seqn <= main_genericstandalone_rtio_core_sed_record142_rec_seqn;
			main_genericstandalone_rtio_core_sed_record158_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record142_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record158_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record142_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record142_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record142_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_address <= main_genericstandalone_rtio_core_sed_record142_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_data <= main_genericstandalone_rtio_core_sed_record142_rec_payload_data;
		end else begin
			main_genericstandalone_rtio_core_sed_record157_rec_valid <= main_genericstandalone_rtio_core_sed_record142_rec_valid;
			main_genericstandalone_rtio_core_sed_record157_rec_seqn <= main_genericstandalone_rtio_core_sed_record142_rec_seqn;
			main_genericstandalone_rtio_core_sed_record157_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record142_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record157_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record142_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record142_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record142_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_address <= main_genericstandalone_rtio_core_sed_record142_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record157_rec_payload_data <= main_genericstandalone_rtio_core_sed_record142_rec_payload_data;
			main_genericstandalone_rtio_core_sed_record158_rec_valid <= main_genericstandalone_rtio_core_sed_record141_rec_valid;
			main_genericstandalone_rtio_core_sed_record158_rec_seqn <= main_genericstandalone_rtio_core_sed_record141_rec_seqn;
			main_genericstandalone_rtio_core_sed_record158_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record141_rec_replace_occured;
			main_genericstandalone_rtio_core_sed_record158_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record141_rec_nondata_replace_occured;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record141_rec_payload_channel;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record141_rec_payload_fine_ts;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_address <= main_genericstandalone_rtio_core_sed_record141_rec_payload_address;
			main_genericstandalone_rtio_core_sed_record158_rec_payload_data <= main_genericstandalone_rtio_core_sed_record141_rec_payload_data;
		end
	end
	main_genericstandalone_rtio_core_sed_record144_rec_valid <= main_genericstandalone_rtio_core_sed_record128_rec_valid;
	main_genericstandalone_rtio_core_sed_record144_rec_seqn <= main_genericstandalone_rtio_core_sed_record128_rec_seqn;
	main_genericstandalone_rtio_core_sed_record144_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record128_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record144_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record128_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record144_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record128_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record144_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record128_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record144_rec_payload_address <= main_genericstandalone_rtio_core_sed_record128_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record144_rec_payload_data <= main_genericstandalone_rtio_core_sed_record128_rec_payload_data;
	main_genericstandalone_rtio_core_sed_record159_rec_valid <= main_genericstandalone_rtio_core_sed_record143_rec_valid;
	main_genericstandalone_rtio_core_sed_record159_rec_seqn <= main_genericstandalone_rtio_core_sed_record143_rec_seqn;
	main_genericstandalone_rtio_core_sed_record159_rec_replace_occured <= main_genericstandalone_rtio_core_sed_record143_rec_replace_occured;
	main_genericstandalone_rtio_core_sed_record159_rec_nondata_replace_occured <= main_genericstandalone_rtio_core_sed_record143_rec_nondata_replace_occured;
	main_genericstandalone_rtio_core_sed_record159_rec_payload_channel <= main_genericstandalone_rtio_core_sed_record143_rec_payload_channel;
	main_genericstandalone_rtio_core_sed_record159_rec_payload_fine_ts <= main_genericstandalone_rtio_core_sed_record143_rec_payload_fine_ts;
	main_genericstandalone_rtio_core_sed_record159_rec_payload_address <= main_genericstandalone_rtio_core_sed_record143_rec_payload_address;
	main_genericstandalone_rtio_core_sed_record159_rec_payload_data <= main_genericstandalone_rtio_core_sed_record143_rec_payload_data;
	if ((main_genericstandalone_rtio_core_inputcollector_selected0 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow0 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger0) begin
		main_genericstandalone_rtio_core_inputcollector_overflow0 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_inputcollector_selected1 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow1 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger1) begin
		main_genericstandalone_rtio_core_inputcollector_overflow1 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_inputcollector_selected2 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow2 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger2) begin
		main_genericstandalone_rtio_core_inputcollector_overflow2 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_inputcollector_selected3 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow3 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger3) begin
		main_genericstandalone_rtio_core_inputcollector_overflow3 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_inputcollector_selected4 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow4 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger4) begin
		main_genericstandalone_rtio_core_inputcollector_overflow4 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_inputcollector_selected5 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow5 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger5) begin
		main_genericstandalone_rtio_core_inputcollector_overflow5 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_inputcollector_selected6 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow6 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger6) begin
		main_genericstandalone_rtio_core_inputcollector_overflow6 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_inputcollector_selected7 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow7 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger7) begin
		main_genericstandalone_rtio_core_inputcollector_overflow7 <= 1'd1;
	end
	if ((main_genericstandalone_rtio_core_inputcollector_selected8 & main_genericstandalone_rtio_core_inputcollector_i_ack)) begin
		main_genericstandalone_rtio_core_inputcollector_overflow8 <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_inputcollector_overflow_trigger8) begin
		main_genericstandalone_rtio_core_inputcollector_overflow8 <= 1'd1;
	end
	main_genericstandalone_rtio_core_inputcollector_i_ack <= 1'd0;
	if (main_genericstandalone_rtio_core_inputcollector_i_ack) begin
		main_genericstandalone_rtio_core_cri_i_status <= {1'd0, main_genericstandalone_rtio_core_inputcollector_i_status_raw[1], (~main_genericstandalone_rtio_core_inputcollector_i_status_raw[0])};
		main_genericstandalone_rtio_core_cri_i_data <= builder_sync_t_rhs_self1;
		main_genericstandalone_rtio_core_cri_i_timestamp <= builder_sync_t_rhs_self2;
	end
	if (((main_genericstandalone_full_ts >= main_genericstandalone_rtio_core_inputcollector_input_timeout) | (main_genericstandalone_rtio_core_inputcollector_i_status_raw != 1'd0))) begin
		if (main_genericstandalone_rtio_core_inputcollector_input_pending) begin
			main_genericstandalone_rtio_core_inputcollector_i_ack <= 1'd1;
		end
		main_genericstandalone_rtio_core_inputcollector_input_pending <= 1'd0;
	end
	if ((main_genericstandalone_rtio_core_cri_cmd == 2'd2)) begin
		main_genericstandalone_rtio_core_inputcollector_input_timeout <= main_genericstandalone_rtio_core_cri_i_timeout;
		main_genericstandalone_rtio_core_inputcollector_input_pending <= 1'd1;
		main_genericstandalone_rtio_core_cri_i_status <= 3'd4;
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_syncfifo0_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_syncfifo1_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_syncfifo2_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_syncfifo3_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_syncfifo4_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_syncfifo5_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_syncfifo6_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_syncfifo7_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_re) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_re) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_replace))) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_produce <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_do_read) begin
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_consume <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_we & main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_syncfifo8_writable) & (~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_replace))) begin
		if ((~main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_do_read)) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_do_read) begin
			main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 <= (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 - 1'd1);
		end
	end
	if (main_genericstandalone_rtio_core_o_collision_sync_i) begin
		main_genericstandalone_rtio_core_o_collision_sync_blind <= 1'd1;
	end
	if (main_genericstandalone_rtio_core_o_collision_sync_ps_ack_o) begin
		main_genericstandalone_rtio_core_o_collision_sync_blind <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_o_collision_sync_ps_i) begin
		main_genericstandalone_rtio_core_o_collision_sync_bxfer_data <= main_genericstandalone_rtio_core_o_collision_sync_data_i;
	end
	if (main_genericstandalone_rtio_core_o_collision_sync_ps_i) begin
		main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_i <= (~main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_i);
	end
	main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_o_r <= main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_o;
	if (main_genericstandalone_rtio_core_o_busy_sync_i) begin
		main_genericstandalone_rtio_core_o_busy_sync_blind <= 1'd1;
	end
	if (main_genericstandalone_rtio_core_o_busy_sync_ps_ack_o) begin
		main_genericstandalone_rtio_core_o_busy_sync_blind <= 1'd0;
	end
	if (main_genericstandalone_rtio_core_o_busy_sync_ps_i) begin
		main_genericstandalone_rtio_core_o_busy_sync_bxfer_data <= main_genericstandalone_rtio_core_o_busy_sync_data_i;
	end
	if (main_genericstandalone_rtio_core_o_busy_sync_ps_i) begin
		main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_i <= (~main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_i);
	end
	main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_o_r <= main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_o;
	main_genericstandalone_mon_bussynchronizer20_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer20_pong_o) begin
		main_genericstandalone_mon_bussynchronizer20_ibuffer <= main_genericstandalone_mon_bussynchronizer20_i;
	end
	if (main_genericstandalone_mon_bussynchronizer20_ping_i) begin
		main_genericstandalone_mon_bussynchronizer20_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer20_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer20_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer20_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer20_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer20_done)) begin
			main_genericstandalone_mon_bussynchronizer20_count <= (main_genericstandalone_mon_bussynchronizer20_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer20_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer21_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer21_pong_o) begin
		main_genericstandalone_mon_bussynchronizer21_ibuffer <= main_genericstandalone_mon_bussynchronizer21_i;
	end
	if (main_genericstandalone_mon_bussynchronizer21_ping_i) begin
		main_genericstandalone_mon_bussynchronizer21_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer21_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer21_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer21_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer21_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer21_done)) begin
			main_genericstandalone_mon_bussynchronizer21_count <= (main_genericstandalone_mon_bussynchronizer21_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer21_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer22_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer22_pong_o) begin
		main_genericstandalone_mon_bussynchronizer22_ibuffer <= main_genericstandalone_mon_bussynchronizer22_i;
	end
	if (main_genericstandalone_mon_bussynchronizer22_ping_i) begin
		main_genericstandalone_mon_bussynchronizer22_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer22_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer22_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer22_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer22_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer22_done)) begin
			main_genericstandalone_mon_bussynchronizer22_count <= (main_genericstandalone_mon_bussynchronizer22_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer22_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer23_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer23_pong_o) begin
		main_genericstandalone_mon_bussynchronizer23_ibuffer <= main_genericstandalone_mon_bussynchronizer23_i;
	end
	if (main_genericstandalone_mon_bussynchronizer23_ping_i) begin
		main_genericstandalone_mon_bussynchronizer23_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer23_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer23_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer23_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer23_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer23_done)) begin
			main_genericstandalone_mon_bussynchronizer23_count <= (main_genericstandalone_mon_bussynchronizer23_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer23_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer29_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer29_pong_o) begin
		main_genericstandalone_mon_bussynchronizer29_ibuffer <= main_genericstandalone_mon_bussynchronizer29_i;
	end
	if (main_genericstandalone_mon_bussynchronizer29_ping_i) begin
		main_genericstandalone_mon_bussynchronizer29_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer29_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer29_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer29_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer29_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer29_done)) begin
			main_genericstandalone_mon_bussynchronizer29_count <= (main_genericstandalone_mon_bussynchronizer29_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer29_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer30_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer30_pong_o) begin
		main_genericstandalone_mon_bussynchronizer30_ibuffer <= main_genericstandalone_mon_bussynchronizer30_i;
	end
	if (main_genericstandalone_mon_bussynchronizer30_ping_i) begin
		main_genericstandalone_mon_bussynchronizer30_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer30_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer30_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer30_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer30_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer30_done)) begin
			main_genericstandalone_mon_bussynchronizer30_count <= (main_genericstandalone_mon_bussynchronizer30_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer30_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer31_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer31_pong_o) begin
		main_genericstandalone_mon_bussynchronizer31_ibuffer <= main_genericstandalone_mon_bussynchronizer31_i;
	end
	if (main_genericstandalone_mon_bussynchronizer31_ping_i) begin
		main_genericstandalone_mon_bussynchronizer31_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer31_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer31_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer31_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer31_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer31_done)) begin
			main_genericstandalone_mon_bussynchronizer31_count <= (main_genericstandalone_mon_bussynchronizer31_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer31_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer32_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer32_pong_o) begin
		main_genericstandalone_mon_bussynchronizer32_ibuffer <= main_genericstandalone_mon_bussynchronizer32_i;
	end
	if (main_genericstandalone_mon_bussynchronizer32_ping_i) begin
		main_genericstandalone_mon_bussynchronizer32_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer32_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer32_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer32_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer32_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer32_done)) begin
			main_genericstandalone_mon_bussynchronizer32_count <= (main_genericstandalone_mon_bussynchronizer32_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer32_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer39_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer39_pong_o) begin
		main_genericstandalone_mon_bussynchronizer39_ibuffer <= main_genericstandalone_mon_bussynchronizer39_i;
	end
	if (main_genericstandalone_mon_bussynchronizer39_ping_i) begin
		main_genericstandalone_mon_bussynchronizer39_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer39_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer39_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer39_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer39_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer39_done)) begin
			main_genericstandalone_mon_bussynchronizer39_count <= (main_genericstandalone_mon_bussynchronizer39_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer39_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer40_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer40_pong_o) begin
		main_genericstandalone_mon_bussynchronizer40_ibuffer <= main_genericstandalone_mon_bussynchronizer40_i;
	end
	if (main_genericstandalone_mon_bussynchronizer40_ping_i) begin
		main_genericstandalone_mon_bussynchronizer40_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer40_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer40_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer40_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer40_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer40_done)) begin
			main_genericstandalone_mon_bussynchronizer40_count <= (main_genericstandalone_mon_bussynchronizer40_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer40_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer41_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer41_pong_o) begin
		main_genericstandalone_mon_bussynchronizer41_ibuffer <= main_genericstandalone_mon_bussynchronizer41_i;
	end
	if (main_genericstandalone_mon_bussynchronizer41_ping_i) begin
		main_genericstandalone_mon_bussynchronizer41_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer41_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer41_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer41_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer41_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer41_done)) begin
			main_genericstandalone_mon_bussynchronizer41_count <= (main_genericstandalone_mon_bussynchronizer41_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer41_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer42_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer42_pong_o) begin
		main_genericstandalone_mon_bussynchronizer42_ibuffer <= main_genericstandalone_mon_bussynchronizer42_i;
	end
	if (main_genericstandalone_mon_bussynchronizer42_ping_i) begin
		main_genericstandalone_mon_bussynchronizer42_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer42_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer42_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer42_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer42_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer42_done)) begin
			main_genericstandalone_mon_bussynchronizer42_count <= (main_genericstandalone_mon_bussynchronizer42_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer42_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer43_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer43_pong_o) begin
		main_genericstandalone_mon_bussynchronizer43_ibuffer <= main_genericstandalone_mon_bussynchronizer43_i;
	end
	if (main_genericstandalone_mon_bussynchronizer43_ping_i) begin
		main_genericstandalone_mon_bussynchronizer43_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer43_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer43_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer43_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer43_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer43_done)) begin
			main_genericstandalone_mon_bussynchronizer43_count <= (main_genericstandalone_mon_bussynchronizer43_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer43_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer44_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer44_pong_o) begin
		main_genericstandalone_mon_bussynchronizer44_ibuffer <= main_genericstandalone_mon_bussynchronizer44_i;
	end
	if (main_genericstandalone_mon_bussynchronizer44_ping_i) begin
		main_genericstandalone_mon_bussynchronizer44_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer44_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer44_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer44_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer44_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer44_done)) begin
			main_genericstandalone_mon_bussynchronizer44_count <= (main_genericstandalone_mon_bussynchronizer44_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer44_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer45_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer45_pong_o) begin
		main_genericstandalone_mon_bussynchronizer45_ibuffer <= main_genericstandalone_mon_bussynchronizer45_i;
	end
	if (main_genericstandalone_mon_bussynchronizer45_ping_i) begin
		main_genericstandalone_mon_bussynchronizer45_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer45_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer45_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer45_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer45_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer45_done)) begin
			main_genericstandalone_mon_bussynchronizer45_count <= (main_genericstandalone_mon_bussynchronizer45_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer45_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer46_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer46_pong_o) begin
		main_genericstandalone_mon_bussynchronizer46_ibuffer <= main_genericstandalone_mon_bussynchronizer46_i;
	end
	if (main_genericstandalone_mon_bussynchronizer46_ping_i) begin
		main_genericstandalone_mon_bussynchronizer46_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer46_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer46_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer46_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer46_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer46_done)) begin
			main_genericstandalone_mon_bussynchronizer46_count <= (main_genericstandalone_mon_bussynchronizer46_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer46_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer47_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer47_pong_o) begin
		main_genericstandalone_mon_bussynchronizer47_ibuffer <= main_genericstandalone_mon_bussynchronizer47_i;
	end
	if (main_genericstandalone_mon_bussynchronizer47_ping_i) begin
		main_genericstandalone_mon_bussynchronizer47_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer47_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer47_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer47_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer47_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer47_done)) begin
			main_genericstandalone_mon_bussynchronizer47_count <= (main_genericstandalone_mon_bussynchronizer47_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer47_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer48_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer48_pong_o) begin
		main_genericstandalone_mon_bussynchronizer48_ibuffer <= main_genericstandalone_mon_bussynchronizer48_i;
	end
	if (main_genericstandalone_mon_bussynchronizer48_ping_i) begin
		main_genericstandalone_mon_bussynchronizer48_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer48_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer48_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer48_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer48_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer48_done)) begin
			main_genericstandalone_mon_bussynchronizer48_count <= (main_genericstandalone_mon_bussynchronizer48_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer48_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer49_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer49_pong_o) begin
		main_genericstandalone_mon_bussynchronizer49_ibuffer <= main_genericstandalone_mon_bussynchronizer49_i;
	end
	if (main_genericstandalone_mon_bussynchronizer49_ping_i) begin
		main_genericstandalone_mon_bussynchronizer49_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer49_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer49_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer49_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer49_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer49_done)) begin
			main_genericstandalone_mon_bussynchronizer49_count <= (main_genericstandalone_mon_bussynchronizer49_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer49_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer50_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer50_pong_o) begin
		main_genericstandalone_mon_bussynchronizer50_ibuffer <= main_genericstandalone_mon_bussynchronizer50_i;
	end
	if (main_genericstandalone_mon_bussynchronizer50_ping_i) begin
		main_genericstandalone_mon_bussynchronizer50_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer50_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer50_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer50_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer50_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer50_done)) begin
			main_genericstandalone_mon_bussynchronizer50_count <= (main_genericstandalone_mon_bussynchronizer50_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer50_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer51_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer51_pong_o) begin
		main_genericstandalone_mon_bussynchronizer51_ibuffer <= main_genericstandalone_mon_bussynchronizer51_i;
	end
	if (main_genericstandalone_mon_bussynchronizer51_ping_i) begin
		main_genericstandalone_mon_bussynchronizer51_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer51_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer51_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer51_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer51_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer51_done)) begin
			main_genericstandalone_mon_bussynchronizer51_count <= (main_genericstandalone_mon_bussynchronizer51_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer51_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer52_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer52_pong_o) begin
		main_genericstandalone_mon_bussynchronizer52_ibuffer <= main_genericstandalone_mon_bussynchronizer52_i;
	end
	if (main_genericstandalone_mon_bussynchronizer52_ping_i) begin
		main_genericstandalone_mon_bussynchronizer52_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer52_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer52_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer52_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer52_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer52_done)) begin
			main_genericstandalone_mon_bussynchronizer52_count <= (main_genericstandalone_mon_bussynchronizer52_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer52_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer53_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer53_pong_o) begin
		main_genericstandalone_mon_bussynchronizer53_ibuffer <= main_genericstandalone_mon_bussynchronizer53_i;
	end
	if (main_genericstandalone_mon_bussynchronizer53_ping_i) begin
		main_genericstandalone_mon_bussynchronizer53_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer53_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer53_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer53_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer53_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer53_done)) begin
			main_genericstandalone_mon_bussynchronizer53_count <= (main_genericstandalone_mon_bussynchronizer53_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer53_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer54_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer54_pong_o) begin
		main_genericstandalone_mon_bussynchronizer54_ibuffer <= main_genericstandalone_mon_bussynchronizer54_i;
	end
	if (main_genericstandalone_mon_bussynchronizer54_ping_i) begin
		main_genericstandalone_mon_bussynchronizer54_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer54_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer54_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer54_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer54_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer54_done)) begin
			main_genericstandalone_mon_bussynchronizer54_count <= (main_genericstandalone_mon_bussynchronizer54_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer54_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer55_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer55_pong_o) begin
		main_genericstandalone_mon_bussynchronizer55_ibuffer <= main_genericstandalone_mon_bussynchronizer55_i;
	end
	if (main_genericstandalone_mon_bussynchronizer55_ping_i) begin
		main_genericstandalone_mon_bussynchronizer55_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer55_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer55_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer55_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer55_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer55_done)) begin
			main_genericstandalone_mon_bussynchronizer55_count <= (main_genericstandalone_mon_bussynchronizer55_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer55_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer56_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer56_pong_o) begin
		main_genericstandalone_mon_bussynchronizer56_ibuffer <= main_genericstandalone_mon_bussynchronizer56_i;
	end
	if (main_genericstandalone_mon_bussynchronizer56_ping_i) begin
		main_genericstandalone_mon_bussynchronizer56_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer56_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer56_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer56_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer56_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer56_done)) begin
			main_genericstandalone_mon_bussynchronizer56_count <= (main_genericstandalone_mon_bussynchronizer56_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer56_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer57_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer57_pong_o) begin
		main_genericstandalone_mon_bussynchronizer57_ibuffer <= main_genericstandalone_mon_bussynchronizer57_i;
	end
	if (main_genericstandalone_mon_bussynchronizer57_ping_i) begin
		main_genericstandalone_mon_bussynchronizer57_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer57_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer57_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer57_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer57_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer57_done)) begin
			main_genericstandalone_mon_bussynchronizer57_count <= (main_genericstandalone_mon_bussynchronizer57_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer57_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer58_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer58_pong_o) begin
		main_genericstandalone_mon_bussynchronizer58_ibuffer <= main_genericstandalone_mon_bussynchronizer58_i;
	end
	if (main_genericstandalone_mon_bussynchronizer58_ping_i) begin
		main_genericstandalone_mon_bussynchronizer58_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer58_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer58_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer58_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer58_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer58_done)) begin
			main_genericstandalone_mon_bussynchronizer58_count <= (main_genericstandalone_mon_bussynchronizer58_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer58_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer59_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer59_pong_o) begin
		main_genericstandalone_mon_bussynchronizer59_ibuffer <= main_genericstandalone_mon_bussynchronizer59_i;
	end
	if (main_genericstandalone_mon_bussynchronizer59_ping_i) begin
		main_genericstandalone_mon_bussynchronizer59_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer59_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer59_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer59_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer59_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer59_done)) begin
			main_genericstandalone_mon_bussynchronizer59_count <= (main_genericstandalone_mon_bussynchronizer59_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer59_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer60_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer60_pong_o) begin
		main_genericstandalone_mon_bussynchronizer60_ibuffer <= main_genericstandalone_mon_bussynchronizer60_i;
	end
	if (main_genericstandalone_mon_bussynchronizer60_ping_i) begin
		main_genericstandalone_mon_bussynchronizer60_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer60_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer60_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer60_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer60_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer60_done)) begin
			main_genericstandalone_mon_bussynchronizer60_count <= (main_genericstandalone_mon_bussynchronizer60_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer60_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer61_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer61_pong_o) begin
		main_genericstandalone_mon_bussynchronizer61_ibuffer <= main_genericstandalone_mon_bussynchronizer61_i;
	end
	if (main_genericstandalone_mon_bussynchronizer61_ping_i) begin
		main_genericstandalone_mon_bussynchronizer61_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer61_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer61_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer61_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer61_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer61_done)) begin
			main_genericstandalone_mon_bussynchronizer61_count <= (main_genericstandalone_mon_bussynchronizer61_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer61_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer62_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer62_pong_o) begin
		main_genericstandalone_mon_bussynchronizer62_ibuffer <= main_genericstandalone_mon_bussynchronizer62_i;
	end
	if (main_genericstandalone_mon_bussynchronizer62_ping_i) begin
		main_genericstandalone_mon_bussynchronizer62_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer62_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer62_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer62_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer62_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer62_done)) begin
			main_genericstandalone_mon_bussynchronizer62_count <= (main_genericstandalone_mon_bussynchronizer62_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer62_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer63_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer63_pong_o) begin
		main_genericstandalone_mon_bussynchronizer63_ibuffer <= main_genericstandalone_mon_bussynchronizer63_i;
	end
	if (main_genericstandalone_mon_bussynchronizer63_ping_i) begin
		main_genericstandalone_mon_bussynchronizer63_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer63_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer63_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer63_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer63_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer63_done)) begin
			main_genericstandalone_mon_bussynchronizer63_count <= (main_genericstandalone_mon_bussynchronizer63_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer63_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer64_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer64_pong_o) begin
		main_genericstandalone_mon_bussynchronizer64_ibuffer <= main_genericstandalone_mon_bussynchronizer64_i;
	end
	if (main_genericstandalone_mon_bussynchronizer64_ping_i) begin
		main_genericstandalone_mon_bussynchronizer64_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer64_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer64_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer64_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer64_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer64_done)) begin
			main_genericstandalone_mon_bussynchronizer64_count <= (main_genericstandalone_mon_bussynchronizer64_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer64_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer65_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer65_pong_o) begin
		main_genericstandalone_mon_bussynchronizer65_ibuffer <= main_genericstandalone_mon_bussynchronizer65_i;
	end
	if (main_genericstandalone_mon_bussynchronizer65_ping_i) begin
		main_genericstandalone_mon_bussynchronizer65_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer65_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer65_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer65_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer65_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer65_done)) begin
			main_genericstandalone_mon_bussynchronizer65_count <= (main_genericstandalone_mon_bussynchronizer65_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer65_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer66_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer66_pong_o) begin
		main_genericstandalone_mon_bussynchronizer66_ibuffer <= main_genericstandalone_mon_bussynchronizer66_i;
	end
	if (main_genericstandalone_mon_bussynchronizer66_ping_i) begin
		main_genericstandalone_mon_bussynchronizer66_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer66_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer66_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer66_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer66_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer66_done)) begin
			main_genericstandalone_mon_bussynchronizer66_count <= (main_genericstandalone_mon_bussynchronizer66_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer66_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer67_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer67_pong_o) begin
		main_genericstandalone_mon_bussynchronizer67_ibuffer <= main_genericstandalone_mon_bussynchronizer67_i;
	end
	if (main_genericstandalone_mon_bussynchronizer67_ping_i) begin
		main_genericstandalone_mon_bussynchronizer67_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer67_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer67_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer67_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer67_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer67_done)) begin
			main_genericstandalone_mon_bussynchronizer67_count <= (main_genericstandalone_mon_bussynchronizer67_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer67_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer68_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer68_pong_o) begin
		main_genericstandalone_mon_bussynchronizer68_ibuffer <= main_genericstandalone_mon_bussynchronizer68_i;
	end
	if (main_genericstandalone_mon_bussynchronizer68_ping_i) begin
		main_genericstandalone_mon_bussynchronizer68_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer68_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer68_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer68_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer68_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer68_done)) begin
			main_genericstandalone_mon_bussynchronizer68_count <= (main_genericstandalone_mon_bussynchronizer68_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer68_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer69_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer69_pong_o) begin
		main_genericstandalone_mon_bussynchronizer69_ibuffer <= main_genericstandalone_mon_bussynchronizer69_i;
	end
	if (main_genericstandalone_mon_bussynchronizer69_ping_i) begin
		main_genericstandalone_mon_bussynchronizer69_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer69_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer69_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer69_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer69_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer69_done)) begin
			main_genericstandalone_mon_bussynchronizer69_count <= (main_genericstandalone_mon_bussynchronizer69_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer69_count <= 8'd128;
	end
	main_genericstandalone_mon_bussynchronizer70_starter <= 1'd0;
	if (main_genericstandalone_mon_bussynchronizer70_pong_o) begin
		main_genericstandalone_mon_bussynchronizer70_ibuffer <= main_genericstandalone_mon_bussynchronizer70_i;
	end
	if (main_genericstandalone_mon_bussynchronizer70_ping_i) begin
		main_genericstandalone_mon_bussynchronizer70_ping_toggle_i <= (~main_genericstandalone_mon_bussynchronizer70_ping_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer70_pong_toggle_o_r <= main_genericstandalone_mon_bussynchronizer70_pong_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer70_wait) begin
		if ((~main_genericstandalone_mon_bussynchronizer70_done)) begin
			main_genericstandalone_mon_bussynchronizer70_count <= (main_genericstandalone_mon_bussynchronizer70_count - 1'd1);
		end
	end else begin
		main_genericstandalone_mon_bussynchronizer70_count <= 8'd128;
	end
	if (rio_rst) begin
		main_inout_8x0_inout_8x0_ointerface0_stb <= 1'd0;
		main_inout_8x0_inout_8x0_sensitivity <= 2'd0;
		main_inout_8x0_inout_8x0_sample <= 1'd0;
		main_inout_8x1_inout_8x1_ointerface1_stb <= 1'd0;
		main_inout_8x1_inout_8x1_sensitivity <= 2'd0;
		main_inout_8x1_inout_8x1_sample <= 1'd0;
		main_inout_8x2_inout_8x2_ointerface2_stb <= 1'd0;
		main_inout_8x2_inout_8x2_sensitivity <= 2'd0;
		main_inout_8x2_inout_8x2_sample <= 1'd0;
		main_inout_8x3_inout_8x3_ointerface3_stb <= 1'd0;
		main_inout_8x3_inout_8x3_sensitivity <= 2'd0;
		main_inout_8x3_inout_8x3_sample <= 1'd0;
		main_output_8x0_stb0 <= 1'd0;
		main_output_8x1_stb0 <= 1'd0;
		main_output_8x2_stb <= 1'd0;
		main_output_8x3_stb <= 1'd0;
		main_output_8x4_stb <= 1'd0;
		main_output_8x5_stb <= 1'd0;
		main_output_8x6_stb <= 1'd0;
		main_output_8x7_stb <= 1'd0;
		main_output_8x8_stb <= 1'd0;
		main_output_8x9_stb <= 1'd0;
		main_output_8x10_stb <= 1'd0;
		main_output_8x11_stb <= 1'd0;
		main_spimaster0_ointerface0_stb0 <= 1'd0;
		main_output_8x0_stb1 <= 1'd0;
		main_urukulmonitor0_cs <= 8'd0;
		main_urukulmonitor0_data_length <= 8'd0;
		main_urukulmonitor0_flags <= 8'd0;
		main_output_8x12_stb <= 1'd0;
		main_output_8x13_stb <= 1'd0;
		main_output_8x14_stb <= 1'd0;
		main_output_8x15_stb <= 1'd0;
		main_spimaster1_ointerface1_stb0 <= 1'd0;
		main_output_8x1_stb1 <= 1'd0;
		main_urukulmonitor1_cs <= 8'd0;
		main_urukulmonitor1_data_length <= 8'd0;
		main_urukulmonitor1_flags <= 8'd0;
		main_output_8x16_stb <= 1'd0;
		main_output_8x17_stb <= 1'd0;
		main_output_8x18_stb <= 1'd0;
		main_output_8x19_stb <= 1'd0;
		main_spimaster0_ointerface0_stb1 <= 1'd0;
		main_spimaster1_ointerface1_stb1 <= 1'd0;
		main_output_8x20_stb <= 1'd0;
		main_spimaster2_ointerface2_stb <= 1'd0;
		main_ldac_phy_stb <= 1'd0;
		main_clr_phy_stb <= 1'd0;
		main_output0_stb <= 1'd0;
		main_output1_stb <= 1'd0;
		main_output2_stb <= 1'd0;
		main_stb <= 1'd0;
		main_genericstandalone_rtio_core_cri_i_status <= 4'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_sequence_error <= 1'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_o_status_underflow <= 1'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_current_lane <= 4'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_coarse_timestamp <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps0 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps1 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps2 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps3 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps4 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps5 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps6 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps7 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps8 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps9 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps10 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps11 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps12 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps13 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps14 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_last_lane_coarse_timestamps15 <= 61'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_seqn <= 13'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_quash <= 1'd0;
		main_genericstandalone_rtio_core_sed_lane_dist_force_laneB <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered0_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered1_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered2_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered3_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered4_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered5_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered6_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered7_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered8_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered9_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered10_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered11_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered12_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered13_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered14_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_readable <= 1'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_level0 <= 8'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_produce <= 7'd0;
		main_genericstandalone_rtio_core_sed_syncfifobuffered15_consume <= 7'd0;
		main_genericstandalone_rtio_core_sed_gates_record16_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record17_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record18_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record19_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record20_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record21_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record22_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record23_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record24_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record25_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record26_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record27_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record28_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record29_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record30_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_gates_record31_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_collision <= 1'd0;
		main_genericstandalone_rtio_core_sed_busy <= 1'd0;
		main_genericstandalone_rtio_core_sed_record0_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record1_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record2_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record3_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record4_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record5_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record6_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record7_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record8_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record9_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record10_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record11_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record12_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record13_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record14_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record15_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record16_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record17_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record18_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record19_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record20_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record21_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record22_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record23_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record24_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record25_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record26_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record27_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record28_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record29_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record30_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record31_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record32_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record33_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record34_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record35_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record36_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record37_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record38_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record39_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record40_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record41_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record42_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record43_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record44_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record45_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record46_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record47_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record48_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record49_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record50_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record51_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record52_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record53_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record54_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record55_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record56_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record57_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record58_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record59_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record60_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record61_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record62_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record63_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record64_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record65_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record66_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record67_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record68_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record69_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record70_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record71_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record72_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record73_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record74_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record75_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record76_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record77_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record78_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record79_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record80_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record81_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record82_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record83_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record84_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record85_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record86_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record87_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record88_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record89_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record90_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record91_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record92_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record93_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record94_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record95_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record96_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record97_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record98_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record99_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record100_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record101_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record102_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record103_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record104_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record105_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record106_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record107_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record108_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record109_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record110_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record111_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record112_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record113_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record114_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record115_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record116_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record117_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record118_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record119_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record120_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record121_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record122_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record123_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record124_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record125_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record126_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record127_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record128_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record129_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record130_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record131_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record132_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record133_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record134_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record135_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record136_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record137_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record138_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record139_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record140_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record141_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record142_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record143_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record144_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record145_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record146_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record147_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record148_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record149_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record150_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record151_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record152_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record153_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record154_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record155_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record156_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record157_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record158_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record159_rec_valid <= 1'd0;
		main_genericstandalone_rtio_core_sed_record0_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record1_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record2_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record3_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record4_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record5_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record6_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record7_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record8_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record9_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record10_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record11_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record12_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record13_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record14_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_record15_valid1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r0 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r0 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r2 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r2 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r3 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r3 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r4 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r4 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r5 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r5 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r6 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r6 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r7 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r7 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r8 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r8 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r9 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r9 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r10 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r10 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r11 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r11 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r12 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r12 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r13 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r13 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r14 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r14 <= 1'd0;
		main_genericstandalone_rtio_core_sed_replace_occured_r15 <= 1'd0;
		main_genericstandalone_rtio_core_sed_nondata_replace_occured_r15 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r0 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r1 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r2 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r3 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r4 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r5 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r6 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r7 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r8 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r9 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r10 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r11 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r12 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r13 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r14 <= 1'd0;
		main_genericstandalone_rtio_core_sed_stb_r15 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_i_ack <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_level0 <= 7'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_produce <= 6'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_consume <= 6'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow0 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_level0 <= 7'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_produce <= 6'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_consume <= 6'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow1 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_level0 <= 7'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_produce <= 6'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_consume <= 6'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow2 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_level0 <= 7'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_produce <= 6'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_consume <= 6'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow3 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_level0 <= 3'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_produce <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_consume <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow4 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_level0 <= 3'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_produce <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_consume <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow5 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_level0 <= 3'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_produce <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_consume <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow6 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_level0 <= 3'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_produce <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_consume <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow7 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_readable <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_level0 <= 3'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_produce <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_consume <= 2'd0;
		main_genericstandalone_rtio_core_inputcollector_overflow8 <= 1'd0;
		main_genericstandalone_rtio_core_inputcollector_input_pending <= 1'd0;
		main_genericstandalone_rtio_core_o_collision_sync_blind <= 1'd0;
		main_genericstandalone_rtio_core_o_busy_sync_blind <= 1'd0;
		main_genericstandalone_mon_bussynchronizer20_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer20_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer21_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer21_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer22_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer22_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer23_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer23_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer29_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer29_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer30_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer30_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer31_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer31_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer32_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer32_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer39_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer39_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer40_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer40_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer41_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer41_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer42_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer42_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer43_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer43_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer44_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer44_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer45_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer45_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer46_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer46_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer47_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer47_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer48_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer48_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer49_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer49_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer50_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer50_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer51_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer51_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer52_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer52_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer53_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer53_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer54_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer54_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer55_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer55_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer56_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer56_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer57_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer57_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer58_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer58_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer59_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer59_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer60_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer60_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer61_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer61_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer62_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer62_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer63_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer63_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer64_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer64_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer65_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer65_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer66_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer66_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer67_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer67_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer68_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer68_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer69_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer69_count <= 8'd128;
		main_genericstandalone_mon_bussynchronizer70_starter <= 1'd1;
		main_genericstandalone_mon_bussynchronizer70_count <= 8'd128;
	end
	builder_xilinxmultiregimpl210 <= main_genericstandalone_rtio_core_storage;
	builder_xilinxmultiregimpl211 <= builder_xilinxmultiregimpl210;
	builder_xilinxmultiregimpl230 <= main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_i;
	builder_xilinxmultiregimpl231 <= builder_xilinxmultiregimpl230;
	builder_xilinxmultiregimpl260 <= main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_i;
	builder_xilinxmultiregimpl261 <= builder_xilinxmultiregimpl260;
	builder_xilinxmultiregimpl490 <= main_genericstandalone_mon_bussynchronizer20_pong_toggle_i;
	builder_xilinxmultiregimpl491 <= builder_xilinxmultiregimpl490;
	builder_xilinxmultiregimpl520 <= main_genericstandalone_mon_bussynchronizer21_pong_toggle_i;
	builder_xilinxmultiregimpl521 <= builder_xilinxmultiregimpl520;
	builder_xilinxmultiregimpl550 <= main_genericstandalone_mon_bussynchronizer22_pong_toggle_i;
	builder_xilinxmultiregimpl551 <= builder_xilinxmultiregimpl550;
	builder_xilinxmultiregimpl580 <= main_genericstandalone_mon_bussynchronizer23_pong_toggle_i;
	builder_xilinxmultiregimpl581 <= builder_xilinxmultiregimpl580;
	builder_xilinxmultiregimpl660 <= main_genericstandalone_mon_bussynchronizer29_pong_toggle_i;
	builder_xilinxmultiregimpl661 <= builder_xilinxmultiregimpl660;
	builder_xilinxmultiregimpl690 <= main_genericstandalone_mon_bussynchronizer30_pong_toggle_i;
	builder_xilinxmultiregimpl691 <= builder_xilinxmultiregimpl690;
	builder_xilinxmultiregimpl720 <= main_genericstandalone_mon_bussynchronizer31_pong_toggle_i;
	builder_xilinxmultiregimpl721 <= builder_xilinxmultiregimpl720;
	builder_xilinxmultiregimpl750 <= main_genericstandalone_mon_bussynchronizer32_pong_toggle_i;
	builder_xilinxmultiregimpl751 <= builder_xilinxmultiregimpl750;
	builder_xilinxmultiregimpl840 <= main_genericstandalone_mon_bussynchronizer39_pong_toggle_i;
	builder_xilinxmultiregimpl841 <= builder_xilinxmultiregimpl840;
	builder_xilinxmultiregimpl870 <= main_genericstandalone_mon_bussynchronizer40_pong_toggle_i;
	builder_xilinxmultiregimpl871 <= builder_xilinxmultiregimpl870;
	builder_xilinxmultiregimpl900 <= main_genericstandalone_mon_bussynchronizer41_pong_toggle_i;
	builder_xilinxmultiregimpl901 <= builder_xilinxmultiregimpl900;
	builder_xilinxmultiregimpl930 <= main_genericstandalone_mon_bussynchronizer42_pong_toggle_i;
	builder_xilinxmultiregimpl931 <= builder_xilinxmultiregimpl930;
	builder_xilinxmultiregimpl960 <= main_genericstandalone_mon_bussynchronizer43_pong_toggle_i;
	builder_xilinxmultiregimpl961 <= builder_xilinxmultiregimpl960;
	builder_xilinxmultiregimpl990 <= main_genericstandalone_mon_bussynchronizer44_pong_toggle_i;
	builder_xilinxmultiregimpl991 <= builder_xilinxmultiregimpl990;
	builder_xilinxmultiregimpl1020 <= main_genericstandalone_mon_bussynchronizer45_pong_toggle_i;
	builder_xilinxmultiregimpl1021 <= builder_xilinxmultiregimpl1020;
	builder_xilinxmultiregimpl1050 <= main_genericstandalone_mon_bussynchronizer46_pong_toggle_i;
	builder_xilinxmultiregimpl1051 <= builder_xilinxmultiregimpl1050;
	builder_xilinxmultiregimpl1080 <= main_genericstandalone_mon_bussynchronizer47_pong_toggle_i;
	builder_xilinxmultiregimpl1081 <= builder_xilinxmultiregimpl1080;
	builder_xilinxmultiregimpl1110 <= main_genericstandalone_mon_bussynchronizer48_pong_toggle_i;
	builder_xilinxmultiregimpl1111 <= builder_xilinxmultiregimpl1110;
	builder_xilinxmultiregimpl1140 <= main_genericstandalone_mon_bussynchronizer49_pong_toggle_i;
	builder_xilinxmultiregimpl1141 <= builder_xilinxmultiregimpl1140;
	builder_xilinxmultiregimpl1170 <= main_genericstandalone_mon_bussynchronizer50_pong_toggle_i;
	builder_xilinxmultiregimpl1171 <= builder_xilinxmultiregimpl1170;
	builder_xilinxmultiregimpl1200 <= main_genericstandalone_mon_bussynchronizer51_pong_toggle_i;
	builder_xilinxmultiregimpl1201 <= builder_xilinxmultiregimpl1200;
	builder_xilinxmultiregimpl1230 <= main_genericstandalone_mon_bussynchronizer52_pong_toggle_i;
	builder_xilinxmultiregimpl1231 <= builder_xilinxmultiregimpl1230;
	builder_xilinxmultiregimpl1260 <= main_genericstandalone_mon_bussynchronizer53_pong_toggle_i;
	builder_xilinxmultiregimpl1261 <= builder_xilinxmultiregimpl1260;
	builder_xilinxmultiregimpl1290 <= main_genericstandalone_mon_bussynchronizer54_pong_toggle_i;
	builder_xilinxmultiregimpl1291 <= builder_xilinxmultiregimpl1290;
	builder_xilinxmultiregimpl1320 <= main_genericstandalone_mon_bussynchronizer55_pong_toggle_i;
	builder_xilinxmultiregimpl1321 <= builder_xilinxmultiregimpl1320;
	builder_xilinxmultiregimpl1350 <= main_genericstandalone_mon_bussynchronizer56_pong_toggle_i;
	builder_xilinxmultiregimpl1351 <= builder_xilinxmultiregimpl1350;
	builder_xilinxmultiregimpl1380 <= main_genericstandalone_mon_bussynchronizer57_pong_toggle_i;
	builder_xilinxmultiregimpl1381 <= builder_xilinxmultiregimpl1380;
	builder_xilinxmultiregimpl1410 <= main_genericstandalone_mon_bussynchronizer58_pong_toggle_i;
	builder_xilinxmultiregimpl1411 <= builder_xilinxmultiregimpl1410;
	builder_xilinxmultiregimpl1440 <= main_genericstandalone_mon_bussynchronizer59_pong_toggle_i;
	builder_xilinxmultiregimpl1441 <= builder_xilinxmultiregimpl1440;
	builder_xilinxmultiregimpl1470 <= main_genericstandalone_mon_bussynchronizer60_pong_toggle_i;
	builder_xilinxmultiregimpl1471 <= builder_xilinxmultiregimpl1470;
	builder_xilinxmultiregimpl1500 <= main_genericstandalone_mon_bussynchronizer61_pong_toggle_i;
	builder_xilinxmultiregimpl1501 <= builder_xilinxmultiregimpl1500;
	builder_xilinxmultiregimpl1530 <= main_genericstandalone_mon_bussynchronizer62_pong_toggle_i;
	builder_xilinxmultiregimpl1531 <= builder_xilinxmultiregimpl1530;
	builder_xilinxmultiregimpl1560 <= main_genericstandalone_mon_bussynchronizer63_pong_toggle_i;
	builder_xilinxmultiregimpl1561 <= builder_xilinxmultiregimpl1560;
	builder_xilinxmultiregimpl1590 <= main_genericstandalone_mon_bussynchronizer64_pong_toggle_i;
	builder_xilinxmultiregimpl1591 <= builder_xilinxmultiregimpl1590;
	builder_xilinxmultiregimpl1620 <= main_genericstandalone_mon_bussynchronizer65_pong_toggle_i;
	builder_xilinxmultiregimpl1621 <= builder_xilinxmultiregimpl1620;
	builder_xilinxmultiregimpl1650 <= main_genericstandalone_mon_bussynchronizer66_pong_toggle_i;
	builder_xilinxmultiregimpl1651 <= builder_xilinxmultiregimpl1650;
	builder_xilinxmultiregimpl1680 <= main_genericstandalone_mon_bussynchronizer67_pong_toggle_i;
	builder_xilinxmultiregimpl1681 <= builder_xilinxmultiregimpl1680;
	builder_xilinxmultiregimpl1710 <= main_genericstandalone_mon_bussynchronizer68_pong_toggle_i;
	builder_xilinxmultiregimpl1711 <= builder_xilinxmultiregimpl1710;
	builder_xilinxmultiregimpl1740 <= main_genericstandalone_mon_bussynchronizer69_pong_toggle_i;
	builder_xilinxmultiregimpl1741 <= builder_xilinxmultiregimpl1740;
	builder_xilinxmultiregimpl1770 <= main_genericstandalone_mon_bussynchronizer70_pong_toggle_i;
	builder_xilinxmultiregimpl1771 <= builder_xilinxmultiregimpl1770;
	builder_xilinxmultiregimpl1840 <= main_genericstandalone_inj_o_sys0;
	builder_xilinxmultiregimpl1841 <= builder_xilinxmultiregimpl1840;
	builder_xilinxmultiregimpl1850 <= main_genericstandalone_inj_o_sys1;
	builder_xilinxmultiregimpl1851 <= builder_xilinxmultiregimpl1850;
	builder_xilinxmultiregimpl1860 <= main_genericstandalone_inj_o_sys2;
	builder_xilinxmultiregimpl1861 <= builder_xilinxmultiregimpl1860;
	builder_xilinxmultiregimpl1870 <= main_genericstandalone_inj_o_sys3;
	builder_xilinxmultiregimpl1871 <= builder_xilinxmultiregimpl1870;
	builder_xilinxmultiregimpl1880 <= main_genericstandalone_inj_o_sys4;
	builder_xilinxmultiregimpl1881 <= builder_xilinxmultiregimpl1880;
	builder_xilinxmultiregimpl1890 <= main_genericstandalone_inj_o_sys5;
	builder_xilinxmultiregimpl1891 <= builder_xilinxmultiregimpl1890;
	builder_xilinxmultiregimpl1900 <= main_genericstandalone_inj_o_sys6;
	builder_xilinxmultiregimpl1901 <= builder_xilinxmultiregimpl1900;
	builder_xilinxmultiregimpl1910 <= main_genericstandalone_inj_o_sys7;
	builder_xilinxmultiregimpl1911 <= builder_xilinxmultiregimpl1910;
	builder_xilinxmultiregimpl1920 <= main_genericstandalone_inj_o_sys8;
	builder_xilinxmultiregimpl1921 <= builder_xilinxmultiregimpl1920;
	builder_xilinxmultiregimpl1930 <= main_genericstandalone_inj_o_sys9;
	builder_xilinxmultiregimpl1931 <= builder_xilinxmultiregimpl1930;
	builder_xilinxmultiregimpl1940 <= main_genericstandalone_inj_o_sys10;
	builder_xilinxmultiregimpl1941 <= builder_xilinxmultiregimpl1940;
	builder_xilinxmultiregimpl1950 <= main_genericstandalone_inj_o_sys11;
	builder_xilinxmultiregimpl1951 <= builder_xilinxmultiregimpl1950;
	builder_xilinxmultiregimpl1960 <= main_genericstandalone_inj_o_sys12;
	builder_xilinxmultiregimpl1961 <= builder_xilinxmultiregimpl1960;
	builder_xilinxmultiregimpl1970 <= main_genericstandalone_inj_o_sys13;
	builder_xilinxmultiregimpl1971 <= builder_xilinxmultiregimpl1970;
	builder_xilinxmultiregimpl1980 <= main_genericstandalone_inj_o_sys14;
	builder_xilinxmultiregimpl1981 <= builder_xilinxmultiregimpl1980;
	builder_xilinxmultiregimpl1990 <= main_genericstandalone_inj_o_sys15;
	builder_xilinxmultiregimpl1991 <= builder_xilinxmultiregimpl1990;
	builder_xilinxmultiregimpl2000 <= main_genericstandalone_inj_o_sys16;
	builder_xilinxmultiregimpl2001 <= builder_xilinxmultiregimpl2000;
	builder_xilinxmultiregimpl2010 <= main_genericstandalone_inj_o_sys17;
	builder_xilinxmultiregimpl2011 <= builder_xilinxmultiregimpl2010;
	builder_xilinxmultiregimpl2020 <= main_genericstandalone_inj_o_sys18;
	builder_xilinxmultiregimpl2021 <= builder_xilinxmultiregimpl2020;
	builder_xilinxmultiregimpl2030 <= main_genericstandalone_inj_o_sys19;
	builder_xilinxmultiregimpl2031 <= builder_xilinxmultiregimpl2030;
	builder_xilinxmultiregimpl2040 <= main_genericstandalone_inj_o_sys20;
	builder_xilinxmultiregimpl2041 <= builder_xilinxmultiregimpl2040;
	builder_xilinxmultiregimpl2050 <= main_genericstandalone_inj_o_sys21;
	builder_xilinxmultiregimpl2051 <= builder_xilinxmultiregimpl2050;
	builder_xilinxmultiregimpl2060 <= main_genericstandalone_inj_o_sys22;
	builder_xilinxmultiregimpl2061 <= builder_xilinxmultiregimpl2060;
	builder_xilinxmultiregimpl2070 <= main_genericstandalone_inj_o_sys23;
	builder_xilinxmultiregimpl2071 <= builder_xilinxmultiregimpl2070;
	builder_xilinxmultiregimpl2080 <= main_genericstandalone_inj_o_sys24;
	builder_xilinxmultiregimpl2081 <= builder_xilinxmultiregimpl2080;
	builder_xilinxmultiregimpl2090 <= main_genericstandalone_inj_o_sys25;
	builder_xilinxmultiregimpl2091 <= builder_xilinxmultiregimpl2090;
	builder_xilinxmultiregimpl2100 <= main_genericstandalone_inj_o_sys26;
	builder_xilinxmultiregimpl2101 <= builder_xilinxmultiregimpl2100;
	builder_xilinxmultiregimpl2110 <= main_genericstandalone_inj_o_sys27;
	builder_xilinxmultiregimpl2111 <= builder_xilinxmultiregimpl2110;
	builder_xilinxmultiregimpl2120 <= main_genericstandalone_inj_o_sys28;
	builder_xilinxmultiregimpl2121 <= builder_xilinxmultiregimpl2120;
	builder_xilinxmultiregimpl2130 <= main_genericstandalone_inj_o_sys29;
	builder_xilinxmultiregimpl2131 <= builder_xilinxmultiregimpl2130;
	builder_xilinxmultiregimpl2140 <= main_genericstandalone_inj_o_sys30;
	builder_xilinxmultiregimpl2141 <= builder_xilinxmultiregimpl2140;
	builder_xilinxmultiregimpl2150 <= main_genericstandalone_inj_o_sys31;
	builder_xilinxmultiregimpl2151 <= builder_xilinxmultiregimpl2150;
	builder_xilinxmultiregimpl2160 <= main_genericstandalone_inj_o_sys32;
	builder_xilinxmultiregimpl2161 <= builder_xilinxmultiregimpl2160;
	builder_xilinxmultiregimpl2170 <= main_genericstandalone_inj_o_sys33;
	builder_xilinxmultiregimpl2171 <= builder_xilinxmultiregimpl2170;
	builder_xilinxmultiregimpl2180 <= main_genericstandalone_inj_o_sys34;
	builder_xilinxmultiregimpl2181 <= builder_xilinxmultiregimpl2180;
	builder_xilinxmultiregimpl2190 <= main_genericstandalone_inj_o_sys35;
	builder_xilinxmultiregimpl2191 <= builder_xilinxmultiregimpl2190;
	builder_xilinxmultiregimpl2200 <= main_genericstandalone_inj_o_sys36;
	builder_xilinxmultiregimpl2201 <= builder_xilinxmultiregimpl2200;
	builder_xilinxmultiregimpl2210 <= main_genericstandalone_inj_o_sys37;
	builder_xilinxmultiregimpl2211 <= builder_xilinxmultiregimpl2210;
	builder_xilinxmultiregimpl2220 <= main_genericstandalone_inj_o_sys38;
	builder_xilinxmultiregimpl2221 <= builder_xilinxmultiregimpl2220;
	builder_xilinxmultiregimpl2230 <= main_genericstandalone_inj_o_sys39;
	builder_xilinxmultiregimpl2231 <= builder_xilinxmultiregimpl2230;
	builder_xilinxmultiregimpl2240 <= main_genericstandalone_inj_o_sys40;
	builder_xilinxmultiregimpl2241 <= builder_xilinxmultiregimpl2240;
	builder_xilinxmultiregimpl2250 <= main_genericstandalone_inj_o_sys41;
	builder_xilinxmultiregimpl2251 <= builder_xilinxmultiregimpl2250;
	builder_xilinxmultiregimpl2260 <= main_genericstandalone_inj_o_sys42;
	builder_xilinxmultiregimpl2261 <= builder_xilinxmultiregimpl2260;
	builder_xilinxmultiregimpl2270 <= main_genericstandalone_inj_o_sys43;
	builder_xilinxmultiregimpl2271 <= builder_xilinxmultiregimpl2270;
	builder_xilinxmultiregimpl2280 <= main_genericstandalone_inj_o_sys44;
	builder_xilinxmultiregimpl2281 <= builder_xilinxmultiregimpl2280;
	builder_xilinxmultiregimpl2290 <= main_genericstandalone_inj_o_sys45;
	builder_xilinxmultiregimpl2291 <= builder_xilinxmultiregimpl2290;
	builder_xilinxmultiregimpl2300 <= main_genericstandalone_inj_o_sys46;
	builder_xilinxmultiregimpl2301 <= builder_xilinxmultiregimpl2300;
	builder_xilinxmultiregimpl2310 <= main_genericstandalone_inj_o_sys47;
	builder_xilinxmultiregimpl2311 <= builder_xilinxmultiregimpl2310;
	builder_xilinxmultiregimpl2320 <= main_genericstandalone_inj_o_sys48;
	builder_xilinxmultiregimpl2321 <= builder_xilinxmultiregimpl2320;
	builder_xilinxmultiregimpl2330 <= main_genericstandalone_inj_o_sys49;
	builder_xilinxmultiregimpl2331 <= builder_xilinxmultiregimpl2330;
	builder_xilinxmultiregimpl2340 <= main_genericstandalone_inj_o_sys50;
	builder_xilinxmultiregimpl2341 <= builder_xilinxmultiregimpl2340;
	builder_xilinxmultiregimpl2350 <= main_genericstandalone_inj_o_sys51;
	builder_xilinxmultiregimpl2351 <= builder_xilinxmultiregimpl2350;
	builder_xilinxmultiregimpl2360 <= main_genericstandalone_inj_o_sys52;
	builder_xilinxmultiregimpl2361 <= builder_xilinxmultiregimpl2360;
	builder_xilinxmultiregimpl2370 <= main_genericstandalone_inj_o_sys53;
	builder_xilinxmultiregimpl2371 <= builder_xilinxmultiregimpl2370;
	builder_xilinxmultiregimpl2380 <= main_genericstandalone_inj_o_sys54;
	builder_xilinxmultiregimpl2381 <= builder_xilinxmultiregimpl2380;
	builder_xilinxmultiregimpl2390 <= main_genericstandalone_inj_o_sys55;
	builder_xilinxmultiregimpl2391 <= builder_xilinxmultiregimpl2390;
	builder_xilinxmultiregimpl2400 <= main_genericstandalone_inj_o_sys56;
	builder_xilinxmultiregimpl2401 <= builder_xilinxmultiregimpl2400;
	builder_xilinxmultiregimpl2410 <= main_genericstandalone_inj_o_sys57;
	builder_xilinxmultiregimpl2411 <= builder_xilinxmultiregimpl2410;
	builder_xilinxmultiregimpl2420 <= main_genericstandalone_inj_o_sys58;
	builder_xilinxmultiregimpl2421 <= builder_xilinxmultiregimpl2420;
	builder_xilinxmultiregimpl2430 <= main_genericstandalone_inj_o_sys59;
	builder_xilinxmultiregimpl2431 <= builder_xilinxmultiregimpl2430;
	builder_xilinxmultiregimpl2440 <= main_genericstandalone_inj_o_sys60;
	builder_xilinxmultiregimpl2441 <= builder_xilinxmultiregimpl2440;
	builder_xilinxmultiregimpl2450 <= main_genericstandalone_inj_o_sys61;
	builder_xilinxmultiregimpl2451 <= builder_xilinxmultiregimpl2450;
	builder_xilinxmultiregimpl2460 <= main_genericstandalone_inj_o_sys62;
	builder_xilinxmultiregimpl2461 <= builder_xilinxmultiregimpl2460;
	builder_xilinxmultiregimpl2470 <= main_genericstandalone_inj_o_sys63;
	builder_xilinxmultiregimpl2471 <= builder_xilinxmultiregimpl2470;
	builder_xilinxmultiregimpl2480 <= main_genericstandalone_inj_o_sys64;
	builder_xilinxmultiregimpl2481 <= builder_xilinxmultiregimpl2480;
	builder_xilinxmultiregimpl2490 <= main_genericstandalone_inj_o_sys65;
	builder_xilinxmultiregimpl2491 <= builder_xilinxmultiregimpl2490;
	builder_xilinxmultiregimpl2500 <= main_genericstandalone_inj_o_sys66;
	builder_xilinxmultiregimpl2501 <= builder_xilinxmultiregimpl2500;
	builder_xilinxmultiregimpl2510 <= main_genericstandalone_inj_o_sys67;
	builder_xilinxmultiregimpl2511 <= builder_xilinxmultiregimpl2510;
end

always @(posedge rio_phy_clk) begin
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd1))) begin
		main_inout_8x0_inout_8x0_oe_k <= main_inout_8x0_inout_8x0_ointerface0_data[0];
	end
	if (main_inout_8x0_inout_8x0_override_en) begin
		main_inout_8x0_inout_8x0_oe <= main_inout_8x0_inout_8x0_override_oe;
	end else begin
		main_inout_8x0_inout_8x0_oe <= main_inout_8x0_inout_8x0_oe_k;
	end
	main_inout_8x0_inout_8x0_i_d <= main_inout_8x0_serdes_i0[7];
	main_inout_8x0_inout_8x0_iinterface0_data <= main_inout_8x0_serdes_i0[7];
	main_inout_8x0_inout_8x0_iinterface0_fine_ts <= main_inout_8x0_inout_8x0_o;
	main_inout_8x0_inout_8x0_iinterface0_stb <= (main_inout_8x0_inout_8x0_sample | (~main_inout_8x0_inout_8x0_n));
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0))) begin
		main_inout_8x0_inout_8x0_previous_data <= main_inout_8x0_inout_8x0_ointerface0_data[0];
	end
	if (main_inout_8x0_inout_8x0_override_en) begin
		main_inout_8x0_serdes_o0 <= {8{main_inout_8x0_inout_8x0_override_o}};
	end else begin
		if ((((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0)) & (~main_inout_8x0_inout_8x0_previous_data)) & main_inout_8x0_inout_8x0_ointerface0_data[0])) begin
			main_inout_8x0_serdes_o0 <= builder_sync_f_t_self1;
		end else begin
			if ((((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0)) & main_inout_8x0_inout_8x0_previous_data) & (~main_inout_8x0_inout_8x0_ointerface0_data[0]))) begin
				main_inout_8x0_serdes_o0 <= builder_sync_f_t_self2;
			end else begin
				main_inout_8x0_serdes_o0 <= {8{main_inout_8x0_inout_8x0_previous_data}};
			end
		end
	end
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd1))) begin
		main_inout_8x1_inout_8x1_oe_k <= main_inout_8x1_inout_8x1_ointerface1_data[0];
	end
	if (main_inout_8x1_inout_8x1_override_en) begin
		main_inout_8x1_inout_8x1_oe <= main_inout_8x1_inout_8x1_override_oe;
	end else begin
		main_inout_8x1_inout_8x1_oe <= main_inout_8x1_inout_8x1_oe_k;
	end
	main_inout_8x1_inout_8x1_i_d <= main_inout_8x1_serdes_i0[7];
	main_inout_8x1_inout_8x1_iinterface1_data <= main_inout_8x1_serdes_i0[7];
	main_inout_8x1_inout_8x1_iinterface1_fine_ts <= main_inout_8x1_inout_8x1_o;
	main_inout_8x1_inout_8x1_iinterface1_stb <= (main_inout_8x1_inout_8x1_sample | (~main_inout_8x1_inout_8x1_n));
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0))) begin
		main_inout_8x1_inout_8x1_previous_data <= main_inout_8x1_inout_8x1_ointerface1_data[0];
	end
	if (main_inout_8x1_inout_8x1_override_en) begin
		main_inout_8x1_serdes_o0 <= {8{main_inout_8x1_inout_8x1_override_o}};
	end else begin
		if ((((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0)) & (~main_inout_8x1_inout_8x1_previous_data)) & main_inout_8x1_inout_8x1_ointerface1_data[0])) begin
			main_inout_8x1_serdes_o0 <= builder_sync_f_t_self3;
		end else begin
			if ((((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0)) & main_inout_8x1_inout_8x1_previous_data) & (~main_inout_8x1_inout_8x1_ointerface1_data[0]))) begin
				main_inout_8x1_serdes_o0 <= builder_sync_f_t_self4;
			end else begin
				main_inout_8x1_serdes_o0 <= {8{main_inout_8x1_inout_8x1_previous_data}};
			end
		end
	end
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd1))) begin
		main_inout_8x2_inout_8x2_oe_k <= main_inout_8x2_inout_8x2_ointerface2_data[0];
	end
	if (main_inout_8x2_inout_8x2_override_en) begin
		main_inout_8x2_inout_8x2_oe <= main_inout_8x2_inout_8x2_override_oe;
	end else begin
		main_inout_8x2_inout_8x2_oe <= main_inout_8x2_inout_8x2_oe_k;
	end
	main_inout_8x2_inout_8x2_i_d <= main_inout_8x2_serdes_i0[7];
	main_inout_8x2_inout_8x2_iinterface2_data <= main_inout_8x2_serdes_i0[7];
	main_inout_8x2_inout_8x2_iinterface2_fine_ts <= main_inout_8x2_inout_8x2_o;
	main_inout_8x2_inout_8x2_iinterface2_stb <= (main_inout_8x2_inout_8x2_sample | (~main_inout_8x2_inout_8x2_n));
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0))) begin
		main_inout_8x2_inout_8x2_previous_data <= main_inout_8x2_inout_8x2_ointerface2_data[0];
	end
	if (main_inout_8x2_inout_8x2_override_en) begin
		main_inout_8x2_serdes_o0 <= {8{main_inout_8x2_inout_8x2_override_o}};
	end else begin
		if ((((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0)) & (~main_inout_8x2_inout_8x2_previous_data)) & main_inout_8x2_inout_8x2_ointerface2_data[0])) begin
			main_inout_8x2_serdes_o0 <= builder_sync_f_t_self5;
		end else begin
			if ((((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0)) & main_inout_8x2_inout_8x2_previous_data) & (~main_inout_8x2_inout_8x2_ointerface2_data[0]))) begin
				main_inout_8x2_serdes_o0 <= builder_sync_f_t_self6;
			end else begin
				main_inout_8x2_serdes_o0 <= {8{main_inout_8x2_inout_8x2_previous_data}};
			end
		end
	end
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd1))) begin
		main_inout_8x3_inout_8x3_oe_k <= main_inout_8x3_inout_8x3_ointerface3_data[0];
	end
	if (main_inout_8x3_inout_8x3_override_en) begin
		main_inout_8x3_inout_8x3_oe <= main_inout_8x3_inout_8x3_override_oe;
	end else begin
		main_inout_8x3_inout_8x3_oe <= main_inout_8x3_inout_8x3_oe_k;
	end
	main_inout_8x3_inout_8x3_i_d <= main_inout_8x3_serdes_i0[7];
	main_inout_8x3_inout_8x3_iinterface3_data <= main_inout_8x3_serdes_i0[7];
	main_inout_8x3_inout_8x3_iinterface3_fine_ts <= main_inout_8x3_inout_8x3_o;
	main_inout_8x3_inout_8x3_iinterface3_stb <= (main_inout_8x3_inout_8x3_sample | (~main_inout_8x3_inout_8x3_n));
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0))) begin
		main_inout_8x3_inout_8x3_previous_data <= main_inout_8x3_inout_8x3_ointerface3_data[0];
	end
	if (main_inout_8x3_inout_8x3_override_en) begin
		main_inout_8x3_serdes_o0 <= {8{main_inout_8x3_inout_8x3_override_o}};
	end else begin
		if ((((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0)) & (~main_inout_8x3_inout_8x3_previous_data)) & main_inout_8x3_inout_8x3_ointerface3_data[0])) begin
			main_inout_8x3_serdes_o0 <= builder_sync_f_t_self7;
		end else begin
			if ((((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0)) & main_inout_8x3_inout_8x3_previous_data) & (~main_inout_8x3_inout_8x3_ointerface3_data[0]))) begin
				main_inout_8x3_serdes_o0 <= builder_sync_f_t_self8;
			end else begin
				main_inout_8x3_serdes_o0 <= {8{main_inout_8x3_inout_8x3_previous_data}};
			end
		end
	end
	if (main_output_8x0_stb0) begin
		main_output_8x0_previous_data0 <= main_output_8x0_data0;
	end
	if (main_output_8x0_override_en0) begin
		main_output_8x0_o0 <= {8{main_output_8x0_override_o0}};
	end else begin
		if (((main_output_8x0_stb0 & (~main_output_8x0_previous_data0)) & main_output_8x0_data0)) begin
			main_output_8x0_o0 <= builder_sync_f_t_self9;
		end else begin
			if (((main_output_8x0_stb0 & main_output_8x0_previous_data0) & (~main_output_8x0_data0))) begin
				main_output_8x0_o0 <= builder_sync_f_t_self10;
			end else begin
				main_output_8x0_o0 <= {8{main_output_8x0_previous_data0}};
			end
		end
	end
	if (main_output_8x1_stb0) begin
		main_output_8x1_previous_data0 <= main_output_8x1_data0;
	end
	if (main_output_8x1_override_en0) begin
		main_output_8x1_o0 <= {8{main_output_8x1_override_o0}};
	end else begin
		if (((main_output_8x1_stb0 & (~main_output_8x1_previous_data0)) & main_output_8x1_data0)) begin
			main_output_8x1_o0 <= builder_sync_f_t_self11;
		end else begin
			if (((main_output_8x1_stb0 & main_output_8x1_previous_data0) & (~main_output_8x1_data0))) begin
				main_output_8x1_o0 <= builder_sync_f_t_self12;
			end else begin
				main_output_8x1_o0 <= {8{main_output_8x1_previous_data0}};
			end
		end
	end
	if (main_output_8x2_stb) begin
		main_output_8x2_previous_data <= main_output_8x2_data;
	end
	if (main_output_8x2_override_en) begin
		main_output_8x2_o <= {8{main_output_8x2_override_o}};
	end else begin
		if (((main_output_8x2_stb & (~main_output_8x2_previous_data)) & main_output_8x2_data)) begin
			main_output_8x2_o <= builder_sync_f_t_self13;
		end else begin
			if (((main_output_8x2_stb & main_output_8x2_previous_data) & (~main_output_8x2_data))) begin
				main_output_8x2_o <= builder_sync_f_t_self14;
			end else begin
				main_output_8x2_o <= {8{main_output_8x2_previous_data}};
			end
		end
	end
	if (main_output_8x3_stb) begin
		main_output_8x3_previous_data <= main_output_8x3_data;
	end
	if (main_output_8x3_override_en) begin
		main_output_8x3_o <= {8{main_output_8x3_override_o}};
	end else begin
		if (((main_output_8x3_stb & (~main_output_8x3_previous_data)) & main_output_8x3_data)) begin
			main_output_8x3_o <= builder_sync_f_t_self15;
		end else begin
			if (((main_output_8x3_stb & main_output_8x3_previous_data) & (~main_output_8x3_data))) begin
				main_output_8x3_o <= builder_sync_f_t_self16;
			end else begin
				main_output_8x3_o <= {8{main_output_8x3_previous_data}};
			end
		end
	end
	if (main_output_8x4_stb) begin
		main_output_8x4_previous_data <= main_output_8x4_data;
	end
	if (main_output_8x4_override_en) begin
		main_output_8x4_o <= {8{main_output_8x4_override_o}};
	end else begin
		if (((main_output_8x4_stb & (~main_output_8x4_previous_data)) & main_output_8x4_data)) begin
			main_output_8x4_o <= builder_sync_f_t_self17;
		end else begin
			if (((main_output_8x4_stb & main_output_8x4_previous_data) & (~main_output_8x4_data))) begin
				main_output_8x4_o <= builder_sync_f_t_self18;
			end else begin
				main_output_8x4_o <= {8{main_output_8x4_previous_data}};
			end
		end
	end
	if (main_output_8x5_stb) begin
		main_output_8x5_previous_data <= main_output_8x5_data;
	end
	if (main_output_8x5_override_en) begin
		main_output_8x5_o <= {8{main_output_8x5_override_o}};
	end else begin
		if (((main_output_8x5_stb & (~main_output_8x5_previous_data)) & main_output_8x5_data)) begin
			main_output_8x5_o <= builder_sync_f_t_self19;
		end else begin
			if (((main_output_8x5_stb & main_output_8x5_previous_data) & (~main_output_8x5_data))) begin
				main_output_8x5_o <= builder_sync_f_t_self20;
			end else begin
				main_output_8x5_o <= {8{main_output_8x5_previous_data}};
			end
		end
	end
	if (main_output_8x6_stb) begin
		main_output_8x6_previous_data <= main_output_8x6_data;
	end
	if (main_output_8x6_override_en) begin
		main_output_8x6_o <= {8{main_output_8x6_override_o}};
	end else begin
		if (((main_output_8x6_stb & (~main_output_8x6_previous_data)) & main_output_8x6_data)) begin
			main_output_8x6_o <= builder_sync_f_t_self21;
		end else begin
			if (((main_output_8x6_stb & main_output_8x6_previous_data) & (~main_output_8x6_data))) begin
				main_output_8x6_o <= builder_sync_f_t_self22;
			end else begin
				main_output_8x6_o <= {8{main_output_8x6_previous_data}};
			end
		end
	end
	if (main_output_8x7_stb) begin
		main_output_8x7_previous_data <= main_output_8x7_data;
	end
	if (main_output_8x7_override_en) begin
		main_output_8x7_o <= {8{main_output_8x7_override_o}};
	end else begin
		if (((main_output_8x7_stb & (~main_output_8x7_previous_data)) & main_output_8x7_data)) begin
			main_output_8x7_o <= builder_sync_f_t_self23;
		end else begin
			if (((main_output_8x7_stb & main_output_8x7_previous_data) & (~main_output_8x7_data))) begin
				main_output_8x7_o <= builder_sync_f_t_self24;
			end else begin
				main_output_8x7_o <= {8{main_output_8x7_previous_data}};
			end
		end
	end
	if (main_output_8x8_stb) begin
		main_output_8x8_previous_data <= main_output_8x8_data;
	end
	if (main_output_8x8_override_en) begin
		main_output_8x8_o <= {8{main_output_8x8_override_o}};
	end else begin
		if (((main_output_8x8_stb & (~main_output_8x8_previous_data)) & main_output_8x8_data)) begin
			main_output_8x8_o <= builder_sync_f_t_self25;
		end else begin
			if (((main_output_8x8_stb & main_output_8x8_previous_data) & (~main_output_8x8_data))) begin
				main_output_8x8_o <= builder_sync_f_t_self26;
			end else begin
				main_output_8x8_o <= {8{main_output_8x8_previous_data}};
			end
		end
	end
	if (main_output_8x9_stb) begin
		main_output_8x9_previous_data <= main_output_8x9_data;
	end
	if (main_output_8x9_override_en) begin
		main_output_8x9_o <= {8{main_output_8x9_override_o}};
	end else begin
		if (((main_output_8x9_stb & (~main_output_8x9_previous_data)) & main_output_8x9_data)) begin
			main_output_8x9_o <= builder_sync_f_t_self27;
		end else begin
			if (((main_output_8x9_stb & main_output_8x9_previous_data) & (~main_output_8x9_data))) begin
				main_output_8x9_o <= builder_sync_f_t_self28;
			end else begin
				main_output_8x9_o <= {8{main_output_8x9_previous_data}};
			end
		end
	end
	if (main_output_8x10_stb) begin
		main_output_8x10_previous_data <= main_output_8x10_data;
	end
	if (main_output_8x10_override_en) begin
		main_output_8x10_o <= {8{main_output_8x10_override_o}};
	end else begin
		if (((main_output_8x10_stb & (~main_output_8x10_previous_data)) & main_output_8x10_data)) begin
			main_output_8x10_o <= builder_sync_f_t_self29;
		end else begin
			if (((main_output_8x10_stb & main_output_8x10_previous_data) & (~main_output_8x10_data))) begin
				main_output_8x10_o <= builder_sync_f_t_self30;
			end else begin
				main_output_8x10_o <= {8{main_output_8x10_previous_data}};
			end
		end
	end
	if (main_output_8x11_stb) begin
		main_output_8x11_previous_data <= main_output_8x11_data;
	end
	if (main_output_8x11_override_en) begin
		main_output_8x11_o <= {8{main_output_8x11_override_o}};
	end else begin
		if (((main_output_8x11_stb & (~main_output_8x11_previous_data)) & main_output_8x11_data)) begin
			main_output_8x11_o <= builder_sync_f_t_self31;
		end else begin
			if (((main_output_8x11_stb & main_output_8x11_previous_data) & (~main_output_8x11_data))) begin
				main_output_8x11_o <= builder_sync_f_t_self32;
			end else begin
				main_output_8x11_o <= {8{main_output_8x11_previous_data}};
			end
		end
	end
	if (main_spimaster0_iinterface0_stb0) begin
		main_spimaster0_read0 <= 1'd0;
	end
	if ((main_spimaster0_ointerface0_stb0 & main_spimaster0_spimachine0_writable0)) begin
		if (main_spimaster0_ointerface0_address0) begin
			{main_spimaster0_config_cs0, main_spimaster0_config_div0, main_spimaster0_config_padding0, main_spimaster0_config_length0, main_spimaster0_config_half_duplex0, main_spimaster0_config_lsb_first0, main_spimaster0_config_clk_phase0, main_spimaster0_config_clk_polarity0, main_spimaster0_config_cs_polarity0, main_spimaster0_config_input0, main_spimaster0_config_end0, main_spimaster0_config_offline0} <= main_spimaster0_ointerface0_data0;
		end else begin
			main_spimaster0_read0 <= main_spimaster0_config_input0;
		end
	end
	if (main_spimaster0_interface_ce0) begin
		main_spimaster0_interface_cs1 <= (({3{main_spimaster0_interface_cs_next0}} & main_spimaster0_interface_cs0) ^ (~main_spimaster0_interface_cs_polarity0));
		main_spimaster0_interface_clk0 <= (main_spimaster0_interface_clk_next0 ^ main_spimaster0_interface_clk_polarity0);
	end
	if (main_spimaster0_interface_sample0) begin
		main_spimaster0_interface_miso_reg0 <= main_spimaster0_interface_miso0;
		main_spimaster0_interface_mosi_reg0 <= main_spimaster0_interface_mosi0;
	end
	if (main_spimaster0_spimachine0_load1) begin
		main_spimaster0_spimachine0_n0 <= main_spimaster0_spimachine0_length0;
		main_spimaster0_spimachine0_end1 <= main_spimaster0_spimachine0_end0;
	end
	if (main_spimaster0_spimachine0_shift0) begin
		main_spimaster0_spimachine0_n0 <= (main_spimaster0_spimachine0_n0 - 1'd1);
	end
	if (main_spimaster0_spimachine0_shift0) begin
		main_spimaster0_spimachine0_sr0 <= main_spimaster0_spimachine0_pdi0;
		main_spimaster0_spimachine0_sdo0 <= (main_spimaster0_spimachine0_lsb_first0 ? main_spimaster0_spimachine0_pdi0[0] : main_spimaster0_spimachine0_pdi0[31]);
	end
	if (main_spimaster0_spimachine0_load1) begin
		main_spimaster0_spimachine0_sr0 <= main_spimaster0_spimachine0_pdo0;
		main_spimaster0_spimachine0_sdo0 <= (main_spimaster0_spimachine0_lsb_first0 ? main_spimaster0_spimachine0_pdo0[0] : main_spimaster0_spimachine0_pdo0[31]);
	end
	if (main_spimaster0_spimachine0_count0) begin
		if (main_spimaster0_spimachine0_cnt_done0) begin
			if (main_spimaster0_spimachine0_do_extend0) begin
				main_spimaster0_spimachine0_do_extend0 <= 1'd0;
			end else begin
				main_spimaster0_spimachine0_cnt0 <= main_spimaster0_spimachine0_div0[7:1];
				main_spimaster0_spimachine0_do_extend0 <= (main_spimaster0_spimachine0_extend0 & main_spimaster0_spimachine0_div0[0]);
			end
		end else begin
			main_spimaster0_spimachine0_cnt0 <= (main_spimaster0_spimachine0_cnt0 - 1'd1);
		end
	end
	builder_spimaster0_state <= builder_spimaster0_next_state;
	if (main_output_8x0_stb1) begin
		main_output_8x0_previous_data1 <= main_output_8x0_data1;
	end
	if (main_output_8x0_override_en1) begin
		main_output_8x0_o1 <= {8{main_output_8x0_override_o1}};
	end else begin
		if (((main_output_8x0_stb1 & (~main_output_8x0_previous_data1)) & main_output_8x0_data1)) begin
			main_output_8x0_o1 <= builder_sync_f_t_self33;
		end else begin
			if (((main_output_8x0_stb1 & main_output_8x0_previous_data1) & (~main_output_8x0_data1))) begin
				main_output_8x0_o1 <= builder_sync_f_t_self34;
			end else begin
				main_output_8x0_o1 <= {8{main_output_8x0_previous_data1}};
			end
		end
	end
	if ((main_urukulmonitor0_ch_sel0 & ((main_output_8x0_stb1 & main_output_8x0_data1) | (((main_urukulmonitor0_cs == 1'd1) & (main_urukulmonitor0_flags & 2'd2)) & (((main_urukulmonitor0_current_data[4] | main_urukulmonitor0_current_data[5]) | main_urukulmonitor0_current_data[6]) | main_urukulmonitor0_current_data[7]))))) begin
		main_urukulmonitor00 <= main_urukulmonitor0_ftw0;
	end
	if ((main_urukulmonitor0_ch_sel1 & ((main_output_8x0_stb1 & main_output_8x0_data1) | (((main_urukulmonitor0_cs == 1'd1) & (main_urukulmonitor0_flags & 2'd2)) & (((main_urukulmonitor0_current_data[4] | main_urukulmonitor0_current_data[5]) | main_urukulmonitor0_current_data[6]) | main_urukulmonitor0_current_data[7]))))) begin
		main_urukulmonitor01 <= main_urukulmonitor0_ftw1;
	end
	if ((main_urukulmonitor0_ch_sel2 & ((main_output_8x0_stb1 & main_output_8x0_data1) | (((main_urukulmonitor0_cs == 1'd1) & (main_urukulmonitor0_flags & 2'd2)) & (((main_urukulmonitor0_current_data[4] | main_urukulmonitor0_current_data[5]) | main_urukulmonitor0_current_data[6]) | main_urukulmonitor0_current_data[7]))))) begin
		main_urukulmonitor02 <= main_urukulmonitor0_ftw2;
	end
	if ((main_urukulmonitor0_ch_sel3 & ((main_output_8x0_stb1 & main_output_8x0_data1) | (((main_urukulmonitor0_cs == 1'd1) & (main_urukulmonitor0_flags & 2'd2)) & (((main_urukulmonitor0_current_data[4] | main_urukulmonitor0_current_data[5]) | main_urukulmonitor0_current_data[6]) | main_urukulmonitor0_current_data[7]))))) begin
		main_urukulmonitor03 <= main_urukulmonitor0_ftw3;
	end
	builder_ad9910monitor0_state <= builder_ad9910monitor0_next_state;
	if (builder_ad9910monitor0_next_value_ce) begin
		main_urukulmonitor0_ftw0[15:0] <= builder_ad9910monitor0_next_value;
	end
	if (main_urukulmonitor0_ftw0_ad9910monitor0_next_value_ce) begin
		main_urukulmonitor0_ftw0 <= main_urukulmonitor0_ftw0_ad9910monitor0_next_value;
	end
	builder_ad9910monitor1_state <= builder_ad9910monitor1_next_state;
	if (builder_ad9910monitor1_next_value_ce) begin
		main_urukulmonitor0_ftw1[15:0] <= builder_ad9910monitor1_next_value;
	end
	if (main_urukulmonitor0_ftw1_ad9910monitor1_next_value_ce) begin
		main_urukulmonitor0_ftw1 <= main_urukulmonitor0_ftw1_ad9910monitor1_next_value;
	end
	builder_ad9910monitor2_state <= builder_ad9910monitor2_next_state;
	if (builder_ad9910monitor2_next_value_ce) begin
		main_urukulmonitor0_ftw2[15:0] <= builder_ad9910monitor2_next_value;
	end
	if (main_urukulmonitor0_ftw2_ad9910monitor2_next_value_ce) begin
		main_urukulmonitor0_ftw2 <= main_urukulmonitor0_ftw2_ad9910monitor2_next_value;
	end
	builder_ad9910monitor3_state <= builder_ad9910monitor3_next_state;
	if (builder_ad9910monitor3_next_value_ce) begin
		main_urukulmonitor0_ftw3[15:0] <= builder_ad9910monitor3_next_value;
	end
	if (main_urukulmonitor0_ftw3_ad9910monitor3_next_value_ce) begin
		main_urukulmonitor0_ftw3 <= main_urukulmonitor0_ftw3_ad9910monitor3_next_value;
	end
	if (main_output_8x12_stb) begin
		main_output_8x12_previous_data <= main_output_8x12_data;
	end
	if (main_output_8x12_override_en) begin
		main_output_8x12_o <= {8{main_output_8x12_override_o}};
	end else begin
		if (((main_output_8x12_stb & (~main_output_8x12_previous_data)) & main_output_8x12_data)) begin
			main_output_8x12_o <= builder_sync_f_t_self35;
		end else begin
			if (((main_output_8x12_stb & main_output_8x12_previous_data) & (~main_output_8x12_data))) begin
				main_output_8x12_o <= builder_sync_f_t_self36;
			end else begin
				main_output_8x12_o <= {8{main_output_8x12_previous_data}};
			end
		end
	end
	if (main_output_8x13_stb) begin
		main_output_8x13_previous_data <= main_output_8x13_data;
	end
	if (main_output_8x13_override_en) begin
		main_output_8x13_o <= {8{main_output_8x13_override_o}};
	end else begin
		if (((main_output_8x13_stb & (~main_output_8x13_previous_data)) & main_output_8x13_data)) begin
			main_output_8x13_o <= builder_sync_f_t_self37;
		end else begin
			if (((main_output_8x13_stb & main_output_8x13_previous_data) & (~main_output_8x13_data))) begin
				main_output_8x13_o <= builder_sync_f_t_self38;
			end else begin
				main_output_8x13_o <= {8{main_output_8x13_previous_data}};
			end
		end
	end
	if (main_output_8x14_stb) begin
		main_output_8x14_previous_data <= main_output_8x14_data;
	end
	if (main_output_8x14_override_en) begin
		main_output_8x14_o <= {8{main_output_8x14_override_o}};
	end else begin
		if (((main_output_8x14_stb & (~main_output_8x14_previous_data)) & main_output_8x14_data)) begin
			main_output_8x14_o <= builder_sync_f_t_self39;
		end else begin
			if (((main_output_8x14_stb & main_output_8x14_previous_data) & (~main_output_8x14_data))) begin
				main_output_8x14_o <= builder_sync_f_t_self40;
			end else begin
				main_output_8x14_o <= {8{main_output_8x14_previous_data}};
			end
		end
	end
	if (main_output_8x15_stb) begin
		main_output_8x15_previous_data <= main_output_8x15_data;
	end
	if (main_output_8x15_override_en) begin
		main_output_8x15_o <= {8{main_output_8x15_override_o}};
	end else begin
		if (((main_output_8x15_stb & (~main_output_8x15_previous_data)) & main_output_8x15_data)) begin
			main_output_8x15_o <= builder_sync_f_t_self41;
		end else begin
			if (((main_output_8x15_stb & main_output_8x15_previous_data) & (~main_output_8x15_data))) begin
				main_output_8x15_o <= builder_sync_f_t_self42;
			end else begin
				main_output_8x15_o <= {8{main_output_8x15_previous_data}};
			end
		end
	end
	if (main_spimaster1_iinterface1_stb0) begin
		main_spimaster1_read0 <= 1'd0;
	end
	if ((main_spimaster1_ointerface1_stb0 & main_spimaster1_spimachine1_writable0)) begin
		if (main_spimaster1_ointerface1_address0) begin
			{main_spimaster1_config_cs0, main_spimaster1_config_div0, main_spimaster1_config_padding0, main_spimaster1_config_length0, main_spimaster1_config_half_duplex0, main_spimaster1_config_lsb_first0, main_spimaster1_config_clk_phase0, main_spimaster1_config_clk_polarity0, main_spimaster1_config_cs_polarity0, main_spimaster1_config_input0, main_spimaster1_config_end0, main_spimaster1_config_offline0} <= main_spimaster1_ointerface1_data0;
		end else begin
			main_spimaster1_read0 <= main_spimaster1_config_input0;
		end
	end
	if (main_spimaster1_interface_ce0) begin
		main_spimaster1_interface_cs1 <= (({3{main_spimaster1_interface_cs_next0}} & main_spimaster1_interface_cs0) ^ (~main_spimaster1_interface_cs_polarity0));
		main_spimaster1_interface_clk0 <= (main_spimaster1_interface_clk_next0 ^ main_spimaster1_interface_clk_polarity0);
	end
	if (main_spimaster1_interface_sample0) begin
		main_spimaster1_interface_miso_reg0 <= main_spimaster1_interface_miso0;
		main_spimaster1_interface_mosi_reg0 <= main_spimaster1_interface_mosi0;
	end
	if (main_spimaster1_spimachine1_load1) begin
		main_spimaster1_spimachine1_n0 <= main_spimaster1_spimachine1_length0;
		main_spimaster1_spimachine1_end1 <= main_spimaster1_spimachine1_end0;
	end
	if (main_spimaster1_spimachine1_shift0) begin
		main_spimaster1_spimachine1_n0 <= (main_spimaster1_spimachine1_n0 - 1'd1);
	end
	if (main_spimaster1_spimachine1_shift0) begin
		main_spimaster1_spimachine1_sr0 <= main_spimaster1_spimachine1_pdi0;
		main_spimaster1_spimachine1_sdo0 <= (main_spimaster1_spimachine1_lsb_first0 ? main_spimaster1_spimachine1_pdi0[0] : main_spimaster1_spimachine1_pdi0[31]);
	end
	if (main_spimaster1_spimachine1_load1) begin
		main_spimaster1_spimachine1_sr0 <= main_spimaster1_spimachine1_pdo0;
		main_spimaster1_spimachine1_sdo0 <= (main_spimaster1_spimachine1_lsb_first0 ? main_spimaster1_spimachine1_pdo0[0] : main_spimaster1_spimachine1_pdo0[31]);
	end
	if (main_spimaster1_spimachine1_count0) begin
		if (main_spimaster1_spimachine1_cnt_done0) begin
			if (main_spimaster1_spimachine1_do_extend0) begin
				main_spimaster1_spimachine1_do_extend0 <= 1'd0;
			end else begin
				main_spimaster1_spimachine1_cnt0 <= main_spimaster1_spimachine1_div0[7:1];
				main_spimaster1_spimachine1_do_extend0 <= (main_spimaster1_spimachine1_extend0 & main_spimaster1_spimachine1_div0[0]);
			end
		end else begin
			main_spimaster1_spimachine1_cnt0 <= (main_spimaster1_spimachine1_cnt0 - 1'd1);
		end
	end
	builder_spimaster1_state <= builder_spimaster1_next_state;
	if (main_output_8x1_stb1) begin
		main_output_8x1_previous_data1 <= main_output_8x1_data1;
	end
	if (main_output_8x1_override_en1) begin
		main_output_8x1_o1 <= {8{main_output_8x1_override_o1}};
	end else begin
		if (((main_output_8x1_stb1 & (~main_output_8x1_previous_data1)) & main_output_8x1_data1)) begin
			main_output_8x1_o1 <= builder_sync_f_t_self43;
		end else begin
			if (((main_output_8x1_stb1 & main_output_8x1_previous_data1) & (~main_output_8x1_data1))) begin
				main_output_8x1_o1 <= builder_sync_f_t_self44;
			end else begin
				main_output_8x1_o1 <= {8{main_output_8x1_previous_data1}};
			end
		end
	end
	if ((main_urukulmonitor1_ch_sel0 & ((main_output_8x1_stb1 & main_output_8x1_data1) | (((main_urukulmonitor1_cs == 1'd1) & (main_urukulmonitor1_flags & 2'd2)) & (((main_urukulmonitor1_current_data[4] | main_urukulmonitor1_current_data[5]) | main_urukulmonitor1_current_data[6]) | main_urukulmonitor1_current_data[7]))))) begin
		main_urukulmonitor10 <= main_urukulmonitor1_ftw0;
	end
	if ((main_urukulmonitor1_ch_sel1 & ((main_output_8x1_stb1 & main_output_8x1_data1) | (((main_urukulmonitor1_cs == 1'd1) & (main_urukulmonitor1_flags & 2'd2)) & (((main_urukulmonitor1_current_data[4] | main_urukulmonitor1_current_data[5]) | main_urukulmonitor1_current_data[6]) | main_urukulmonitor1_current_data[7]))))) begin
		main_urukulmonitor11 <= main_urukulmonitor1_ftw1;
	end
	if ((main_urukulmonitor1_ch_sel2 & ((main_output_8x1_stb1 & main_output_8x1_data1) | (((main_urukulmonitor1_cs == 1'd1) & (main_urukulmonitor1_flags & 2'd2)) & (((main_urukulmonitor1_current_data[4] | main_urukulmonitor1_current_data[5]) | main_urukulmonitor1_current_data[6]) | main_urukulmonitor1_current_data[7]))))) begin
		main_urukulmonitor12 <= main_urukulmonitor1_ftw2;
	end
	if ((main_urukulmonitor1_ch_sel3 & ((main_output_8x1_stb1 & main_output_8x1_data1) | (((main_urukulmonitor1_cs == 1'd1) & (main_urukulmonitor1_flags & 2'd2)) & (((main_urukulmonitor1_current_data[4] | main_urukulmonitor1_current_data[5]) | main_urukulmonitor1_current_data[6]) | main_urukulmonitor1_current_data[7]))))) begin
		main_urukulmonitor13 <= main_urukulmonitor1_ftw3;
	end
	builder_ad9912monitor0_state <= builder_ad9912monitor0_next_state;
	if (builder_ad9912monitor0_t_next_value_ce) begin
		main_urukulmonitor1_ftw0[15:0] <= builder_ad9912monitor0_t_next_value;
	end
	if (builder_ad9912monitor0_f_next_value_ce) begin
		main_urukulmonitor1_ftw0[31:16] <= builder_ad9912monitor0_f_next_value;
	end
	builder_ad9912monitor1_state <= builder_ad9912monitor1_next_state;
	if (builder_ad9912monitor1_t_next_value_ce) begin
		main_urukulmonitor1_ftw1[15:0] <= builder_ad9912monitor1_t_next_value;
	end
	if (builder_ad9912monitor1_f_next_value_ce) begin
		main_urukulmonitor1_ftw1[31:16] <= builder_ad9912monitor1_f_next_value;
	end
	builder_ad9912monitor2_state <= builder_ad9912monitor2_next_state;
	if (builder_ad9912monitor2_t_next_value_ce) begin
		main_urukulmonitor1_ftw2[15:0] <= builder_ad9912monitor2_t_next_value;
	end
	if (builder_ad9912monitor2_f_next_value_ce) begin
		main_urukulmonitor1_ftw2[31:16] <= builder_ad9912monitor2_f_next_value;
	end
	builder_ad9912monitor3_state <= builder_ad9912monitor3_next_state;
	if (builder_ad9912monitor3_t_next_value_ce) begin
		main_urukulmonitor1_ftw3[15:0] <= builder_ad9912monitor3_t_next_value;
	end
	if (builder_ad9912monitor3_f_next_value_ce) begin
		main_urukulmonitor1_ftw3[31:16] <= builder_ad9912monitor3_f_next_value;
	end
	if (main_output_8x16_stb) begin
		main_output_8x16_previous_data <= main_output_8x16_data;
	end
	if (main_output_8x16_override_en) begin
		main_output_8x16_o <= {8{main_output_8x16_override_o}};
	end else begin
		if (((main_output_8x16_stb & (~main_output_8x16_previous_data)) & main_output_8x16_data)) begin
			main_output_8x16_o <= builder_sync_f_t_self45;
		end else begin
			if (((main_output_8x16_stb & main_output_8x16_previous_data) & (~main_output_8x16_data))) begin
				main_output_8x16_o <= builder_sync_f_t_self46;
			end else begin
				main_output_8x16_o <= {8{main_output_8x16_previous_data}};
			end
		end
	end
	if (main_output_8x17_stb) begin
		main_output_8x17_previous_data <= main_output_8x17_data;
	end
	if (main_output_8x17_override_en) begin
		main_output_8x17_o <= {8{main_output_8x17_override_o}};
	end else begin
		if (((main_output_8x17_stb & (~main_output_8x17_previous_data)) & main_output_8x17_data)) begin
			main_output_8x17_o <= builder_sync_f_t_self47;
		end else begin
			if (((main_output_8x17_stb & main_output_8x17_previous_data) & (~main_output_8x17_data))) begin
				main_output_8x17_o <= builder_sync_f_t_self48;
			end else begin
				main_output_8x17_o <= {8{main_output_8x17_previous_data}};
			end
		end
	end
	if (main_output_8x18_stb) begin
		main_output_8x18_previous_data <= main_output_8x18_data;
	end
	if (main_output_8x18_override_en) begin
		main_output_8x18_o <= {8{main_output_8x18_override_o}};
	end else begin
		if (((main_output_8x18_stb & (~main_output_8x18_previous_data)) & main_output_8x18_data)) begin
			main_output_8x18_o <= builder_sync_f_t_self49;
		end else begin
			if (((main_output_8x18_stb & main_output_8x18_previous_data) & (~main_output_8x18_data))) begin
				main_output_8x18_o <= builder_sync_f_t_self50;
			end else begin
				main_output_8x18_o <= {8{main_output_8x18_previous_data}};
			end
		end
	end
	if (main_output_8x19_stb) begin
		main_output_8x19_previous_data <= main_output_8x19_data;
	end
	if (main_output_8x19_override_en) begin
		main_output_8x19_o <= {8{main_output_8x19_override_o}};
	end else begin
		if (((main_output_8x19_stb & (~main_output_8x19_previous_data)) & main_output_8x19_data)) begin
			main_output_8x19_o <= builder_sync_f_t_self51;
		end else begin
			if (((main_output_8x19_stb & main_output_8x19_previous_data) & (~main_output_8x19_data))) begin
				main_output_8x19_o <= builder_sync_f_t_self52;
			end else begin
				main_output_8x19_o <= {8{main_output_8x19_previous_data}};
			end
		end
	end
	if (main_spimaster0_iinterface0_stb1) begin
		main_spimaster0_read1 <= 1'd0;
	end
	if ((main_spimaster0_ointerface0_stb1 & main_spimaster0_spimachine0_writable1)) begin
		if (main_spimaster0_ointerface0_address1) begin
			{main_spimaster0_config_cs1, main_spimaster0_config_div1, main_spimaster0_config_padding1, main_spimaster0_config_length1, main_spimaster0_config_half_duplex1, main_spimaster0_config_lsb_first1, main_spimaster0_config_clk_phase1, main_spimaster0_config_clk_polarity1, main_spimaster0_config_cs_polarity1, main_spimaster0_config_input1, main_spimaster0_config_end1, main_spimaster0_config_offline1} <= main_spimaster0_ointerface0_data1;
		end else begin
			main_spimaster0_read1 <= main_spimaster0_config_input1;
		end
	end
	if (main_spimaster0_interface_ce1) begin
		main_spimaster0_interface_cs3 <= (({1{main_spimaster0_interface_cs_next1}} & main_spimaster0_interface_cs2) ^ (~main_spimaster0_interface_cs_polarity1));
		main_spimaster0_interface_clk1 <= (main_spimaster0_interface_clk_next1 ^ main_spimaster0_interface_clk_polarity1);
	end
	if (main_spimaster0_interface_sample1) begin
		main_spimaster0_interface_miso_reg1 <= main_spimaster0_interface_miso1;
		main_spimaster0_interface_mosi_reg1 <= main_spimaster0_interface_mosi1;
	end
	if (main_spimaster0_spimachine0_load3) begin
		main_spimaster0_spimachine0_n1 <= main_spimaster0_spimachine0_length1;
		main_spimaster0_spimachine0_end3 <= main_spimaster0_spimachine0_end2;
	end
	if (main_spimaster0_spimachine0_shift1) begin
		main_spimaster0_spimachine0_n1 <= (main_spimaster0_spimachine0_n1 - 1'd1);
	end
	if (main_spimaster0_spimachine0_shift1) begin
		main_spimaster0_spimachine0_sr1 <= main_spimaster0_spimachine0_pdi1;
		main_spimaster0_spimachine0_sdo1 <= (main_spimaster0_spimachine0_lsb_first1 ? main_spimaster0_spimachine0_pdi1[0] : main_spimaster0_spimachine0_pdi1[31]);
	end
	if (main_spimaster0_spimachine0_load3) begin
		main_spimaster0_spimachine0_sr1 <= main_spimaster0_spimachine0_pdo1;
		main_spimaster0_spimachine0_sdo1 <= (main_spimaster0_spimachine0_lsb_first1 ? main_spimaster0_spimachine0_pdo1[0] : main_spimaster0_spimachine0_pdo1[31]);
	end
	if (main_spimaster0_spimachine0_count1) begin
		if (main_spimaster0_spimachine0_cnt_done1) begin
			if (main_spimaster0_spimachine0_do_extend1) begin
				main_spimaster0_spimachine0_do_extend1 <= 1'd0;
			end else begin
				main_spimaster0_spimachine0_cnt1 <= main_spimaster0_spimachine0_div1[7:1];
				main_spimaster0_spimachine0_do_extend1 <= (main_spimaster0_spimachine0_extend1 & main_spimaster0_spimachine0_div1[0]);
			end
		end else begin
			main_spimaster0_spimachine0_cnt1 <= (main_spimaster0_spimachine0_cnt1 - 1'd1);
		end
	end
	builder_spimaster2_state <= builder_spimaster2_next_state;
	if (main_spimaster1_iinterface1_stb1) begin
		main_spimaster1_read1 <= 1'd0;
	end
	if ((main_spimaster1_ointerface1_stb1 & main_spimaster1_spimachine1_writable1)) begin
		if (main_spimaster1_ointerface1_address1) begin
			{main_spimaster1_config_cs1, main_spimaster1_config_div1, main_spimaster1_config_padding1, main_spimaster1_config_length1, main_spimaster1_config_half_duplex1, main_spimaster1_config_lsb_first1, main_spimaster1_config_clk_phase1, main_spimaster1_config_clk_polarity1, main_spimaster1_config_cs_polarity1, main_spimaster1_config_input1, main_spimaster1_config_end1, main_spimaster1_config_offline1} <= main_spimaster1_ointerface1_data1;
		end else begin
			main_spimaster1_read1 <= main_spimaster1_config_input1;
		end
	end
	if (main_spimaster1_interface_ce1) begin
		main_spimaster1_interface_cs3 <= (({1{main_spimaster1_interface_cs_next1}} & main_spimaster1_interface_cs2) ^ (~main_spimaster1_interface_cs_polarity1));
		main_spimaster1_interface_clk1 <= (main_spimaster1_interface_clk_next1 ^ main_spimaster1_interface_clk_polarity1);
	end
	if (main_spimaster1_interface_sample1) begin
		main_spimaster1_interface_miso_reg1 <= main_spimaster1_interface_miso1;
		main_spimaster1_interface_mosi_reg1 <= main_spimaster1_interface_mosi1;
	end
	if (main_spimaster1_spimachine1_load3) begin
		main_spimaster1_spimachine1_n1 <= main_spimaster1_spimachine1_length1;
		main_spimaster1_spimachine1_end3 <= main_spimaster1_spimachine1_end2;
	end
	if (main_spimaster1_spimachine1_shift1) begin
		main_spimaster1_spimachine1_n1 <= (main_spimaster1_spimachine1_n1 - 1'd1);
	end
	if (main_spimaster1_spimachine1_shift1) begin
		main_spimaster1_spimachine1_sr1 <= main_spimaster1_spimachine1_pdi1;
		main_spimaster1_spimachine1_sdo1 <= (main_spimaster1_spimachine1_lsb_first1 ? main_spimaster1_spimachine1_pdi1[0] : main_spimaster1_spimachine1_pdi1[31]);
	end
	if (main_spimaster1_spimachine1_load3) begin
		main_spimaster1_spimachine1_sr1 <= main_spimaster1_spimachine1_pdo1;
		main_spimaster1_spimachine1_sdo1 <= (main_spimaster1_spimachine1_lsb_first1 ? main_spimaster1_spimachine1_pdo1[0] : main_spimaster1_spimachine1_pdo1[31]);
	end
	if (main_spimaster1_spimachine1_count1) begin
		if (main_spimaster1_spimachine1_cnt_done1) begin
			if (main_spimaster1_spimachine1_do_extend1) begin
				main_spimaster1_spimachine1_do_extend1 <= 1'd0;
			end else begin
				main_spimaster1_spimachine1_cnt1 <= main_spimaster1_spimachine1_div1[7:1];
				main_spimaster1_spimachine1_do_extend1 <= (main_spimaster1_spimachine1_extend1 & main_spimaster1_spimachine1_div1[0]);
			end
		end else begin
			main_spimaster1_spimachine1_cnt1 <= (main_spimaster1_spimachine1_cnt1 - 1'd1);
		end
	end
	builder_spimaster3_state <= builder_spimaster3_next_state;
	if (main_output_8x20_stb) begin
		main_output_8x20_previous_data <= main_output_8x20_data;
	end
	if (main_output_8x20_override_en) begin
		main_output_8x20_o <= {8{main_output_8x20_override_o}};
	end else begin
		if (((main_output_8x20_stb & (~main_output_8x20_previous_data)) & main_output_8x20_data)) begin
			main_output_8x20_o <= builder_sync_f_t_self53;
		end else begin
			if (((main_output_8x20_stb & main_output_8x20_previous_data) & (~main_output_8x20_data))) begin
				main_output_8x20_o <= builder_sync_f_t_self54;
			end else begin
				main_output_8x20_o <= {8{main_output_8x20_previous_data}};
			end
		end
	end
	if (main_spimaster2_iinterface2_stb) begin
		main_spimaster2_read <= 1'd0;
	end
	if ((main_spimaster2_ointerface2_stb & main_spimaster2_spimachine2_writable)) begin
		if (main_spimaster2_ointerface2_address) begin
			{main_spimaster2_config_cs, main_spimaster2_config_div, main_spimaster2_config_padding, main_spimaster2_config_length, main_spimaster2_config_half_duplex, main_spimaster2_config_lsb_first, main_spimaster2_config_clk_phase, main_spimaster2_config_clk_polarity, main_spimaster2_config_cs_polarity, main_spimaster2_config_input, main_spimaster2_config_end, main_spimaster2_config_offline} <= main_spimaster2_ointerface2_data;
		end else begin
			main_spimaster2_read <= main_spimaster2_config_input;
		end
	end
	if (main_spimaster2_interface_ce) begin
		main_spimaster2_interface_cs1 <= (({2{main_spimaster2_interface_cs_next}} & main_spimaster2_interface_cs0) ^ (~main_spimaster2_interface_cs_polarity));
		main_spimaster2_interface_clk <= (main_spimaster2_interface_clk_next ^ main_spimaster2_interface_clk_polarity);
	end
	if (main_spimaster2_interface_sample) begin
		main_spimaster2_interface_miso_reg <= main_spimaster2_interface_miso;
		main_spimaster2_interface_mosi_reg <= main_spimaster2_interface_mosi;
	end
	if (main_spimaster2_spimachine2_load1) begin
		main_spimaster2_spimachine2_n <= main_spimaster2_spimachine2_length;
		main_spimaster2_spimachine2_end1 <= main_spimaster2_spimachine2_end0;
	end
	if (main_spimaster2_spimachine2_shift) begin
		main_spimaster2_spimachine2_n <= (main_spimaster2_spimachine2_n - 1'd1);
	end
	if (main_spimaster2_spimachine2_shift) begin
		main_spimaster2_spimachine2_sr <= main_spimaster2_spimachine2_pdi;
		main_spimaster2_spimachine2_sdo <= (main_spimaster2_spimachine2_lsb_first ? main_spimaster2_spimachine2_pdi[0] : main_spimaster2_spimachine2_pdi[31]);
	end
	if (main_spimaster2_spimachine2_load1) begin
		main_spimaster2_spimachine2_sr <= main_spimaster2_spimachine2_pdo;
		main_spimaster2_spimachine2_sdo <= (main_spimaster2_spimachine2_lsb_first ? main_spimaster2_spimachine2_pdo[0] : main_spimaster2_spimachine2_pdo[31]);
	end
	if (main_spimaster2_spimachine2_count) begin
		if (main_spimaster2_spimachine2_cnt_done) begin
			if (main_spimaster2_spimachine2_do_extend) begin
				main_spimaster2_spimachine2_do_extend <= 1'd0;
			end else begin
				main_spimaster2_spimachine2_cnt <= main_spimaster2_spimachine2_div[7:1];
				main_spimaster2_spimachine2_do_extend <= (main_spimaster2_spimachine2_extend & main_spimaster2_spimachine2_div[0]);
			end
		end else begin
			main_spimaster2_spimachine2_cnt <= (main_spimaster2_spimachine2_cnt - 1'd1);
		end
	end
	builder_spimaster4_state <= builder_spimaster4_next_state;
	if (main_ldac_phy_stb) begin
		main_ldac_phy_previous_data <= main_ldac_phy_data;
	end
	if (main_ldac_phy_override_en) begin
		main_ldac_phy_o <= {8{main_ldac_phy_override_o}};
	end else begin
		if (((main_ldac_phy_stb & (~main_ldac_phy_previous_data)) & main_ldac_phy_data)) begin
			main_ldac_phy_o <= builder_sync_f_t_self55;
		end else begin
			if (((main_ldac_phy_stb & main_ldac_phy_previous_data) & (~main_ldac_phy_data))) begin
				main_ldac_phy_o <= builder_sync_f_t_self56;
			end else begin
				main_ldac_phy_o <= {8{main_ldac_phy_previous_data}};
			end
		end
	end
	if (main_clr_phy_stb) begin
		main_clr_phy_previous_data <= main_clr_phy_data;
	end
	if (main_clr_phy_override_en) begin
		main_clr_phy_o <= {8{main_clr_phy_override_o}};
	end else begin
		if (((main_clr_phy_stb & (~main_clr_phy_previous_data)) & main_clr_phy_data)) begin
			main_clr_phy_o <= builder_sync_f_t_self57;
		end else begin
			if (((main_clr_phy_stb & main_clr_phy_previous_data) & (~main_clr_phy_data))) begin
				main_clr_phy_o <= builder_sync_f_t_self58;
			end else begin
				main_clr_phy_o <= {8{main_clr_phy_previous_data}};
			end
		end
	end
	if (((main_ldac_phy_stb & 1'd1) & (~main_ldac_phy_data))) begin
		main_ad53xxmonitor0 <= main_ad53xxmonitor32;
		main_ad53xxmonitor1 <= main_ad53xxmonitor33;
		main_ad53xxmonitor2 <= main_ad53xxmonitor34;
		main_ad53xxmonitor3 <= main_ad53xxmonitor35;
		main_ad53xxmonitor4 <= main_ad53xxmonitor36;
		main_ad53xxmonitor5 <= main_ad53xxmonitor37;
		main_ad53xxmonitor6 <= main_ad53xxmonitor38;
		main_ad53xxmonitor7 <= main_ad53xxmonitor39;
		main_ad53xxmonitor8 <= main_ad53xxmonitor40;
		main_ad53xxmonitor9 <= main_ad53xxmonitor41;
		main_ad53xxmonitor10 <= main_ad53xxmonitor42;
		main_ad53xxmonitor11 <= main_ad53xxmonitor43;
		main_ad53xxmonitor12 <= main_ad53xxmonitor44;
		main_ad53xxmonitor13 <= main_ad53xxmonitor45;
		main_ad53xxmonitor14 <= main_ad53xxmonitor46;
		main_ad53xxmonitor15 <= main_ad53xxmonitor47;
		main_ad53xxmonitor16 <= main_ad53xxmonitor48;
		main_ad53xxmonitor17 <= main_ad53xxmonitor49;
		main_ad53xxmonitor18 <= main_ad53xxmonitor50;
		main_ad53xxmonitor19 <= main_ad53xxmonitor51;
		main_ad53xxmonitor20 <= main_ad53xxmonitor52;
		main_ad53xxmonitor21 <= main_ad53xxmonitor53;
		main_ad53xxmonitor22 <= main_ad53xxmonitor54;
		main_ad53xxmonitor23 <= main_ad53xxmonitor55;
		main_ad53xxmonitor24 <= main_ad53xxmonitor56;
		main_ad53xxmonitor25 <= main_ad53xxmonitor57;
		main_ad53xxmonitor26 <= main_ad53xxmonitor58;
		main_ad53xxmonitor27 <= main_ad53xxmonitor59;
		main_ad53xxmonitor28 <= main_ad53xxmonitor60;
		main_ad53xxmonitor29 <= main_ad53xxmonitor61;
		main_ad53xxmonitor30 <= main_ad53xxmonitor62;
		main_ad53xxmonitor31 <= main_ad53xxmonitor63;
	end
	if ((main_spimaster2_ointerface2_stb & (main_spimaster2_ointerface2_address == 1'd1))) begin
		main_ad53xxmonitor_selected <= (main_spimaster2_ointerface2_data[31:24] == 1'd0);
	end
	if ((main_spimaster2_ointerface2_stb & (main_spimaster2_ointerface2_address == 1'd0))) begin
		case (main_spimaster2_ointerface2_data[31:24])
			8'd200: begin
				main_ad53xxmonitor32 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd201: begin
				main_ad53xxmonitor33 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd202: begin
				main_ad53xxmonitor34 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd203: begin
				main_ad53xxmonitor35 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd204: begin
				main_ad53xxmonitor36 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd205: begin
				main_ad53xxmonitor37 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd206: begin
				main_ad53xxmonitor38 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd207: begin
				main_ad53xxmonitor39 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd208: begin
				main_ad53xxmonitor40 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd209: begin
				main_ad53xxmonitor41 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd210: begin
				main_ad53xxmonitor42 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd211: begin
				main_ad53xxmonitor43 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd212: begin
				main_ad53xxmonitor44 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd213: begin
				main_ad53xxmonitor45 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd214: begin
				main_ad53xxmonitor46 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd215: begin
				main_ad53xxmonitor47 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd216: begin
				main_ad53xxmonitor48 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd217: begin
				main_ad53xxmonitor49 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd218: begin
				main_ad53xxmonitor50 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd219: begin
				main_ad53xxmonitor51 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd220: begin
				main_ad53xxmonitor52 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd221: begin
				main_ad53xxmonitor53 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd222: begin
				main_ad53xxmonitor54 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd223: begin
				main_ad53xxmonitor55 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd224: begin
				main_ad53xxmonitor56 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd225: begin
				main_ad53xxmonitor57 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd226: begin
				main_ad53xxmonitor58 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd227: begin
				main_ad53xxmonitor59 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd228: begin
				main_ad53xxmonitor60 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd229: begin
				main_ad53xxmonitor61 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd230: begin
				main_ad53xxmonitor62 <= main_spimaster2_ointerface2_data[23:8];
			end
			8'd231: begin
				main_ad53xxmonitor63 <= main_spimaster2_ointerface2_data[23:8];
			end
		endcase
	end
	if (main_output0_stb) begin
		main_output0_pad_k <= main_output0_data;
	end
	if (main_output0_override_en) begin
		main_output0_pad_o <= main_output0_override_o;
	end else begin
		main_output0_pad_o <= main_output0_pad_k;
	end
	if (main_output1_stb) begin
		main_output1_pad_k <= main_output1_data;
	end
	if (main_output1_override_en) begin
		main_output1_pad_o <= main_output1_override_o;
	end else begin
		main_output1_pad_o <= main_output1_pad_k;
	end
	if (main_output2_stb) begin
		main_output2_pad_k <= main_output2_data;
	end
	if (main_output2_override_en) begin
		main_output2_pad_o <= main_output2_override_o;
	end else begin
		main_output2_pad_o <= main_output2_pad_k;
	end
	if (rio_phy_rst) begin
		main_inout_8x0_serdes_o0 <= 8'd0;
		main_inout_8x0_inout_8x0_iinterface0_stb <= 1'd0;
		main_inout_8x0_inout_8x0_oe <= 1'd0;
		main_inout_8x0_inout_8x0_previous_data <= 1'd0;
		main_inout_8x0_inout_8x0_oe_k <= 1'd0;
		main_inout_8x0_inout_8x0_i_d <= 1'd0;
		main_inout_8x1_serdes_o0 <= 8'd0;
		main_inout_8x1_inout_8x1_iinterface1_stb <= 1'd0;
		main_inout_8x1_inout_8x1_oe <= 1'd0;
		main_inout_8x1_inout_8x1_previous_data <= 1'd0;
		main_inout_8x1_inout_8x1_oe_k <= 1'd0;
		main_inout_8x1_inout_8x1_i_d <= 1'd0;
		main_inout_8x2_serdes_o0 <= 8'd0;
		main_inout_8x2_inout_8x2_iinterface2_stb <= 1'd0;
		main_inout_8x2_inout_8x2_oe <= 1'd0;
		main_inout_8x2_inout_8x2_previous_data <= 1'd0;
		main_inout_8x2_inout_8x2_oe_k <= 1'd0;
		main_inout_8x2_inout_8x2_i_d <= 1'd0;
		main_inout_8x3_serdes_o0 <= 8'd0;
		main_inout_8x3_inout_8x3_iinterface3_stb <= 1'd0;
		main_inout_8x3_inout_8x3_oe <= 1'd0;
		main_inout_8x3_inout_8x3_previous_data <= 1'd0;
		main_inout_8x3_inout_8x3_oe_k <= 1'd0;
		main_inout_8x3_inout_8x3_i_d <= 1'd0;
		main_output_8x0_o0 <= 8'd0;
		main_output_8x0_previous_data0 <= 1'd0;
		main_output_8x1_o0 <= 8'd0;
		main_output_8x1_previous_data0 <= 1'd0;
		main_output_8x2_o <= 8'd0;
		main_output_8x2_previous_data <= 1'd0;
		main_output_8x3_o <= 8'd0;
		main_output_8x3_previous_data <= 1'd0;
		main_output_8x4_o <= 8'd0;
		main_output_8x4_previous_data <= 1'd0;
		main_output_8x5_o <= 8'd0;
		main_output_8x5_previous_data <= 1'd0;
		main_output_8x6_o <= 8'd0;
		main_output_8x6_previous_data <= 1'd0;
		main_output_8x7_o <= 8'd0;
		main_output_8x7_previous_data <= 1'd0;
		main_output_8x8_o <= 8'd0;
		main_output_8x8_previous_data <= 1'd0;
		main_output_8x9_o <= 8'd0;
		main_output_8x9_previous_data <= 1'd0;
		main_output_8x10_o <= 8'd0;
		main_output_8x10_previous_data <= 1'd0;
		main_output_8x11_o <= 8'd0;
		main_output_8x11_previous_data <= 1'd0;
		main_spimaster0_interface_cs1 <= 3'd7;
		main_spimaster0_interface_clk0 <= 1'd0;
		main_spimaster0_spimachine0_cnt0 <= 7'd0;
		main_spimaster0_spimachine0_do_extend0 <= 1'd0;
		main_spimaster0_config_offline0 <= 1'd1;
		main_spimaster0_config_end0 <= 1'd1;
		main_spimaster0_config_input0 <= 1'd0;
		main_spimaster0_config_cs_polarity0 <= 1'd0;
		main_spimaster0_config_clk_polarity0 <= 1'd0;
		main_spimaster0_config_clk_phase0 <= 1'd0;
		main_spimaster0_config_lsb_first0 <= 1'd0;
		main_spimaster0_config_half_duplex0 <= 1'd0;
		main_spimaster0_config_length0 <= 5'd0;
		main_spimaster0_config_padding0 <= 3'd0;
		main_spimaster0_config_div0 <= 8'd0;
		main_spimaster0_config_cs0 <= 8'd0;
		main_spimaster0_read0 <= 1'd0;
		main_output_8x0_o1 <= 8'd0;
		main_output_8x0_previous_data1 <= 1'd0;
		main_urukulmonitor00 <= 32'd0;
		main_urukulmonitor01 <= 32'd0;
		main_urukulmonitor02 <= 32'd0;
		main_urukulmonitor03 <= 32'd0;
		main_output_8x12_o <= 8'd0;
		main_output_8x12_previous_data <= 1'd0;
		main_output_8x13_o <= 8'd0;
		main_output_8x13_previous_data <= 1'd0;
		main_output_8x14_o <= 8'd0;
		main_output_8x14_previous_data <= 1'd0;
		main_output_8x15_o <= 8'd0;
		main_output_8x15_previous_data <= 1'd0;
		main_spimaster1_interface_cs1 <= 3'd7;
		main_spimaster1_interface_clk0 <= 1'd0;
		main_spimaster1_spimachine1_cnt0 <= 7'd0;
		main_spimaster1_spimachine1_do_extend0 <= 1'd0;
		main_spimaster1_config_offline0 <= 1'd1;
		main_spimaster1_config_end0 <= 1'd1;
		main_spimaster1_config_input0 <= 1'd0;
		main_spimaster1_config_cs_polarity0 <= 1'd0;
		main_spimaster1_config_clk_polarity0 <= 1'd0;
		main_spimaster1_config_clk_phase0 <= 1'd0;
		main_spimaster1_config_lsb_first0 <= 1'd0;
		main_spimaster1_config_half_duplex0 <= 1'd0;
		main_spimaster1_config_length0 <= 5'd0;
		main_spimaster1_config_padding0 <= 3'd0;
		main_spimaster1_config_div0 <= 8'd0;
		main_spimaster1_config_cs0 <= 8'd0;
		main_spimaster1_read0 <= 1'd0;
		main_output_8x1_o1 <= 8'd0;
		main_output_8x1_previous_data1 <= 1'd0;
		main_urukulmonitor10 <= 32'd0;
		main_urukulmonitor11 <= 32'd0;
		main_urukulmonitor12 <= 32'd0;
		main_urukulmonitor13 <= 32'd0;
		main_output_8x16_o <= 8'd0;
		main_output_8x16_previous_data <= 1'd0;
		main_output_8x17_o <= 8'd0;
		main_output_8x17_previous_data <= 1'd0;
		main_output_8x18_o <= 8'd0;
		main_output_8x18_previous_data <= 1'd0;
		main_output_8x19_o <= 8'd0;
		main_output_8x19_previous_data <= 1'd0;
		main_spimaster0_interface_cs3 <= 1'd1;
		main_spimaster0_interface_clk1 <= 1'd0;
		main_spimaster0_spimachine0_cnt1 <= 7'd0;
		main_spimaster0_spimachine0_do_extend1 <= 1'd0;
		main_spimaster0_config_offline1 <= 1'd1;
		main_spimaster0_config_end1 <= 1'd1;
		main_spimaster0_config_input1 <= 1'd0;
		main_spimaster0_config_cs_polarity1 <= 1'd0;
		main_spimaster0_config_clk_polarity1 <= 1'd0;
		main_spimaster0_config_clk_phase1 <= 1'd0;
		main_spimaster0_config_lsb_first1 <= 1'd0;
		main_spimaster0_config_half_duplex1 <= 1'd0;
		main_spimaster0_config_length1 <= 5'd0;
		main_spimaster0_config_padding1 <= 3'd0;
		main_spimaster0_config_div1 <= 8'd0;
		main_spimaster0_config_cs1 <= 8'd0;
		main_spimaster0_read1 <= 1'd0;
		main_spimaster1_interface_cs3 <= 1'd1;
		main_spimaster1_interface_clk1 <= 1'd0;
		main_spimaster1_spimachine1_cnt1 <= 7'd0;
		main_spimaster1_spimachine1_do_extend1 <= 1'd0;
		main_spimaster1_config_offline1 <= 1'd1;
		main_spimaster1_config_end1 <= 1'd1;
		main_spimaster1_config_input1 <= 1'd0;
		main_spimaster1_config_cs_polarity1 <= 1'd0;
		main_spimaster1_config_clk_polarity1 <= 1'd0;
		main_spimaster1_config_clk_phase1 <= 1'd0;
		main_spimaster1_config_lsb_first1 <= 1'd0;
		main_spimaster1_config_half_duplex1 <= 1'd0;
		main_spimaster1_config_length1 <= 5'd0;
		main_spimaster1_config_padding1 <= 3'd0;
		main_spimaster1_config_div1 <= 8'd0;
		main_spimaster1_config_cs1 <= 8'd0;
		main_spimaster1_read1 <= 1'd0;
		main_output_8x20_o <= 8'd0;
		main_output_8x20_previous_data <= 1'd0;
		main_spimaster2_interface_cs1 <= 2'd3;
		main_spimaster2_interface_clk <= 1'd0;
		main_spimaster2_spimachine2_cnt <= 7'd0;
		main_spimaster2_spimachine2_do_extend <= 1'd0;
		main_spimaster2_config_offline <= 1'd1;
		main_spimaster2_config_end <= 1'd1;
		main_spimaster2_config_input <= 1'd0;
		main_spimaster2_config_cs_polarity <= 1'd0;
		main_spimaster2_config_clk_polarity <= 1'd0;
		main_spimaster2_config_clk_phase <= 1'd0;
		main_spimaster2_config_lsb_first <= 1'd0;
		main_spimaster2_config_half_duplex <= 1'd0;
		main_spimaster2_config_length <= 5'd0;
		main_spimaster2_config_padding <= 3'd0;
		main_spimaster2_config_div <= 8'd0;
		main_spimaster2_config_cs <= 8'd0;
		main_spimaster2_read <= 1'd0;
		main_ldac_phy_o <= 8'd0;
		main_ldac_phy_previous_data <= 1'd0;
		main_clr_phy_o <= 8'd0;
		main_clr_phy_previous_data <= 1'd0;
		main_ad53xxmonitor0 <= 16'd0;
		main_ad53xxmonitor1 <= 16'd0;
		main_ad53xxmonitor2 <= 16'd0;
		main_ad53xxmonitor3 <= 16'd0;
		main_ad53xxmonitor4 <= 16'd0;
		main_ad53xxmonitor5 <= 16'd0;
		main_ad53xxmonitor6 <= 16'd0;
		main_ad53xxmonitor7 <= 16'd0;
		main_ad53xxmonitor8 <= 16'd0;
		main_ad53xxmonitor9 <= 16'd0;
		main_ad53xxmonitor10 <= 16'd0;
		main_ad53xxmonitor11 <= 16'd0;
		main_ad53xxmonitor12 <= 16'd0;
		main_ad53xxmonitor13 <= 16'd0;
		main_ad53xxmonitor14 <= 16'd0;
		main_ad53xxmonitor15 <= 16'd0;
		main_ad53xxmonitor16 <= 16'd0;
		main_ad53xxmonitor17 <= 16'd0;
		main_ad53xxmonitor18 <= 16'd0;
		main_ad53xxmonitor19 <= 16'd0;
		main_ad53xxmonitor20 <= 16'd0;
		main_ad53xxmonitor21 <= 16'd0;
		main_ad53xxmonitor22 <= 16'd0;
		main_ad53xxmonitor23 <= 16'd0;
		main_ad53xxmonitor24 <= 16'd0;
		main_ad53xxmonitor25 <= 16'd0;
		main_ad53xxmonitor26 <= 16'd0;
		main_ad53xxmonitor27 <= 16'd0;
		main_ad53xxmonitor28 <= 16'd0;
		main_ad53xxmonitor29 <= 16'd0;
		main_ad53xxmonitor30 <= 16'd0;
		main_ad53xxmonitor31 <= 16'd0;
		main_ad53xxmonitor32 <= 16'd0;
		main_ad53xxmonitor33 <= 16'd0;
		main_ad53xxmonitor34 <= 16'd0;
		main_ad53xxmonitor35 <= 16'd0;
		main_ad53xxmonitor36 <= 16'd0;
		main_ad53xxmonitor37 <= 16'd0;
		main_ad53xxmonitor38 <= 16'd0;
		main_ad53xxmonitor39 <= 16'd0;
		main_ad53xxmonitor40 <= 16'd0;
		main_ad53xxmonitor41 <= 16'd0;
		main_ad53xxmonitor42 <= 16'd0;
		main_ad53xxmonitor43 <= 16'd0;
		main_ad53xxmonitor44 <= 16'd0;
		main_ad53xxmonitor45 <= 16'd0;
		main_ad53xxmonitor46 <= 16'd0;
		main_ad53xxmonitor47 <= 16'd0;
		main_ad53xxmonitor48 <= 16'd0;
		main_ad53xxmonitor49 <= 16'd0;
		main_ad53xxmonitor50 <= 16'd0;
		main_ad53xxmonitor51 <= 16'd0;
		main_ad53xxmonitor52 <= 16'd0;
		main_ad53xxmonitor53 <= 16'd0;
		main_ad53xxmonitor54 <= 16'd0;
		main_ad53xxmonitor55 <= 16'd0;
		main_ad53xxmonitor56 <= 16'd0;
		main_ad53xxmonitor57 <= 16'd0;
		main_ad53xxmonitor58 <= 16'd0;
		main_ad53xxmonitor59 <= 16'd0;
		main_ad53xxmonitor60 <= 16'd0;
		main_ad53xxmonitor61 <= 16'd0;
		main_ad53xxmonitor62 <= 16'd0;
		main_ad53xxmonitor63 <= 16'd0;
		main_ad53xxmonitor_selected <= 1'd0;
		main_output0_pad_k <= 1'd0;
		main_output1_pad_k <= 1'd0;
		main_output2_pad_k <= 1'd0;
		builder_spimaster0_state <= 3'd0;
		builder_ad9910monitor0_state <= 1'd0;
		builder_ad9910monitor1_state <= 1'd0;
		builder_ad9910monitor2_state <= 1'd0;
		builder_ad9910monitor3_state <= 1'd0;
		builder_spimaster1_state <= 3'd0;
		builder_ad9912monitor0_state <= 1'd0;
		builder_ad9912monitor1_state <= 1'd0;
		builder_ad9912monitor2_state <= 1'd0;
		builder_ad9912monitor3_state <= 1'd0;
		builder_spimaster2_state <= 3'd0;
		builder_spimaster3_state <= 3'd0;
		builder_spimaster4_state <= 3'd0;
	end
end

always @(posedge sys_clk) begin
	main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack <= 1'd0;
	if (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & (~main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack))) begin
		main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack <= 1'd1;
	end
	main_genericstandalone_genericstandalone_genericstandalone_interface_we <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w <= main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_w;
	main_genericstandalone_genericstandalone_genericstandalone_interface_adr <= main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_adr;
	main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_interface_dat_r;
	if ((main_genericstandalone_genericstandalone_genericstandalone_trigger == 1'd1)) begin
		main_genericstandalone_genericstandalone_genericstandalone_interface_we <= main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_we;
	end
	if ((main_genericstandalone_genericstandalone_genericstandalone_trigger == 2'd2)) begin
		main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack <= 1'd1;
	end
	if ((main_genericstandalone_genericstandalone_genericstandalone_trigger == 2'd3)) begin
		main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack <= 1'd0;
	end
	if ((main_genericstandalone_genericstandalone_genericstandalone_trigger != 1'd0)) begin
		main_genericstandalone_genericstandalone_genericstandalone_trigger <= (main_genericstandalone_genericstandalone_genericstandalone_trigger + 1'd1);
	end else begin
		if ((main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cyc & main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_stb)) begin
			main_genericstandalone_genericstandalone_genericstandalone_trigger <= 1'd1;
		end
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack <= 1'd0;
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_stb & (~main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy)) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack))) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg <= main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_payload_data;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen & main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy)) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount <= (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount + 1'd1);
			if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy <= 1'd0;
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack <= 1'd1;
				end else begin
					serial_tx <= main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg[0];
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg <= {1'd0, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg[7:1]};
				end
			end
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy) begin
		{main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx} <= (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx + main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage);
	end else begin
		{main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx} <= 1'd0;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_r <= main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx;
	if ((~main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy)) begin
		if (((~main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx) & main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_r)) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount <= 1'd0;
		end
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount <= (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount + 1'd1);
			if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount == 1'd0)) begin
				if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx) begin
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy <= 1'd0;
				end
			end else begin
				if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount == 4'd9)) begin
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy <= 1'd0;
					if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx) begin
						main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_payload_data <= main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg;
						main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb <= 1'd1;
					end
				end else begin
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg <= {main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg[7:1]};
				end
			end
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy) begin
		{main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx} <= (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx + main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage);
	end else begin
		{main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx} <= 32'd2147483648;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_clear) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending <= 1'd0;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_tx_old_trigger <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger;
	if (((~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger) & main_genericstandalone_genericstandalone_genericstandalone_uart_tx_old_trigger)) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending <= 1'd1;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending <= 1'd0;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_rx_old_trigger <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger;
	if (((~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger) & main_genericstandalone_genericstandalone_genericstandalone_uart_rx_old_trigger)) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending <= 1'd1;
	end
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we & main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace))) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce + 1'd1);
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume + 1'd1);
	end
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we & main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace))) begin
		if ((~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read)) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level - 1'd1);
		end
	end
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we & main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace))) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce + 1'd1);
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume + 1'd1);
	end
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we & main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace))) begin
		if ((~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read)) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level - 1'd1);
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage) begin
		if ((main_genericstandalone_genericstandalone_genericstandalone_timer0_value == 1'd0)) begin
			main_genericstandalone_genericstandalone_genericstandalone_timer0_value <= main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage;
		end else begin
			main_genericstandalone_genericstandalone_genericstandalone_timer0_value <= (main_genericstandalone_genericstandalone_genericstandalone_timer0_value - 1'd1);
		end
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_value <= main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status <= main_genericstandalone_genericstandalone_genericstandalone_timer0_value;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_clear) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending <= 1'd0;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_old_trigger <= main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger;
	if (((~main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger) & main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_old_trigger)) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending <= 1'd1;
	end
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en0 <= main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_en;
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en1 <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en0;
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en2 <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en1;
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en3 <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en2;
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4 <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en3;
	main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_valid <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4;
	main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_valid <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4;
	main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_valid <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4;
	main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_valid <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4;
	main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en <= {main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en[2:0], main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_en};
	main_genericstandalone_genericstandalone_ddrphy_oe_dqs <= main_genericstandalone_genericstandalone_ddrphy_oe;
	main_genericstandalone_genericstandalone_ddrphy_oe_dq <= main_genericstandalone_genericstandalone_ddrphy_oe;
	if (main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_valid) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_valid) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_valid) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_valid) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_pending_refresh <= 1'd0;
	end
	if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refi_cycles == 1'd0)) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_pending_refresh <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refi_cycles <= 10'd977;
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refi_cycles <= (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refi_cycles - 1'd1);
	end
	if ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_burst)) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col <= {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[6:0], {3{1'd0}}};
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_adr_inc) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col_inc_next;
		end
	end
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_rdvalid_r <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid;
	{main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata} <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_dat_w0;
	{main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_mask, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_mask, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_mask, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_mask} <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_sel0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_dat_w0 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_dat_w1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_sel0 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_sel1;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset0) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset1) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset2) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset3) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset4) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset5) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset6) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset7) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_wait) begin
		if ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_done)) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_count <= (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_count - 1'd1);
		end
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_count <= 3'd4;
	end
	builder_minicon_state <= builder_minicon_next_state;
	main_genericstandalone_genericstandalone_genericstandalone_cache_adr_offset_r <= main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[2:0];
	if (main_genericstandalone_genericstandalone_genericstandalone_cache_adr_inc) begin
		main_genericstandalone_genericstandalone_genericstandalone_cache_adr_offset_r <= main_genericstandalone_genericstandalone_genericstandalone_cache_next_adr_offset;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_cache_word_clr) begin
		main_genericstandalone_genericstandalone_genericstandalone_cache <= 1'd0;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_cache_word_inc) begin
			main_genericstandalone_genericstandalone_genericstandalone_cache <= (main_genericstandalone_genericstandalone_genericstandalone_cache + 1'd1);
		end
	end
	builder_cache_state <= builder_cache_next_state;
	if ((main_genericstandalone_genericstandalone_spiflash_i1 == 1'd0)) begin
		main_genericstandalone_genericstandalone_spiflash_clk <= 1'd1;
		main_genericstandalone_genericstandalone_spiflash_dqi <= main_genericstandalone_genericstandalone_spiflash_i0;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_i1 == 1'd1)) begin
		main_genericstandalone_genericstandalone_spiflash_i1 <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_clk <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_sr <= {main_genericstandalone_genericstandalone_spiflash_sr[61:0], main_genericstandalone_genericstandalone_spiflash_dqi};
	end else begin
		main_genericstandalone_genericstandalone_spiflash_i1 <= (main_genericstandalone_genericstandalone_spiflash_i1 + 1'd1);
	end
	if ((((main_genericstandalone_genericstandalone_spiflash_bus_cyc & main_genericstandalone_genericstandalone_spiflash_bus_stb) & (main_genericstandalone_genericstandalone_spiflash_i1 == 1'd1)) & (main_genericstandalone_genericstandalone_spiflash_trigger == 1'd0))) begin
		main_genericstandalone_genericstandalone_spiflash_dq_oe <= 1'd1;
		main_genericstandalone_genericstandalone_spiflash_cs_n <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_sr[63:48] <= 16'd61423;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_trigger == 5'd16)) begin
		main_genericstandalone_genericstandalone_spiflash_sr[63:40] <= {main_genericstandalone_genericstandalone_spiflash_bus_adr, {3{1'd0}}};
	end
	if ((main_genericstandalone_genericstandalone_spiflash_trigger == 6'd40)) begin
		main_genericstandalone_genericstandalone_spiflash_dq_oe <= 1'd0;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_trigger == 7'd114)) begin
		main_genericstandalone_genericstandalone_spiflash_bus_ack <= 1'd1;
		main_genericstandalone_genericstandalone_spiflash_cs_n <= 1'd1;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_trigger == 7'd115)) begin
		main_genericstandalone_genericstandalone_spiflash_bus_ack <= 1'd0;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_trigger == 7'd117)) begin
	end
	if ((main_genericstandalone_genericstandalone_spiflash_trigger == 7'd117)) begin
		main_genericstandalone_genericstandalone_spiflash_trigger <= 1'd0;
	end else begin
		if ((main_genericstandalone_genericstandalone_spiflash_trigger != 1'd0)) begin
			main_genericstandalone_genericstandalone_spiflash_trigger <= (main_genericstandalone_genericstandalone_spiflash_trigger + 1'd1);
		end else begin
			if (((main_genericstandalone_genericstandalone_spiflash_bus_cyc & main_genericstandalone_genericstandalone_spiflash_bus_stb) & (main_genericstandalone_genericstandalone_spiflash_i1 == 1'd1))) begin
				main_genericstandalone_genericstandalone_spiflash_trigger <= 1'd1;
			end
		end
	end
	if (main_genericstandalone_genericstandalone_icap_counter_rst) begin
		main_genericstandalone_genericstandalone_icap_counter0 <= 1'd1;
	end else begin
		main_genericstandalone_genericstandalone_icap_counter0 <= (main_genericstandalone_genericstandalone_icap_counter0 - 1'd1);
	end
	if (main_genericstandalone_genericstandalone_icap_i) begin
		main_genericstandalone_genericstandalone_icap_toggle_i <= (~main_genericstandalone_genericstandalone_icap_toggle_i);
	end
	main_genericstandalone_tx_mmcm_reset <= (~main_genericstandalone_genericstandalone_qpll_lock);
	if (main_genericstandalone_rx_reset) begin
		main_genericstandalone_cdr_locked <= 1'd0;
		main_genericstandalone_cdr_lock_counter <= 1'd0;
	end else begin
		if ((main_genericstandalone_cdr_lock_counter != 13'd5000)) begin
			main_genericstandalone_cdr_lock_counter <= (main_genericstandalone_cdr_lock_counter + 1'd1);
		end else begin
			main_genericstandalone_cdr_locked <= 1'd1;
		end
	end
	main_genericstandalone_rx_mmcm_reset <= (~main_genericstandalone_cdr_locked);
	main_genericstandalone_tx_init_qpll_reset0 <= main_genericstandalone_tx_init_qpll_reset1;
	main_genericstandalone_tx_init_tx_reset0 <= main_genericstandalone_tx_init_tx_reset1;
	main_genericstandalone_tx_init_tick <= 1'd0;
	if ((main_genericstandalone_tx_init_timer == 6'd63)) begin
		main_genericstandalone_tx_init_tick <= 1'd1;
		main_genericstandalone_tx_init_timer <= 1'd0;
	end else begin
		main_genericstandalone_tx_init_timer <= (main_genericstandalone_tx_init_timer + 1'd1);
	end
	builder_a7_1000basex_gtptxinit_state <= builder_a7_1000basex_gtptxinit_next_state;
	main_genericstandalone_rx_init_rx_reset0 <= main_genericstandalone_rx_init_rx_reset1;
	main_genericstandalone_rx_init_rx_pma_reset_done_r <= main_genericstandalone_rx_init_rx_pma_reset_done1;
	builder_a7_1000basex_gtprxinit_state <= builder_a7_1000basex_gtprxinit_next_state;
	if (main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value_ce) begin
		main_genericstandalone_rx_init_drpvalue <= main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value;
	end
	main_genericstandalone_toggle_o_r <= main_genericstandalone_toggle_o;
	if (main_genericstandalone_ps_preamble_error_o) begin
		main_genericstandalone_preamble_errors_status <= (main_genericstandalone_preamble_errors_status + 1'd1);
	end
	if (main_genericstandalone_ps_crc_error_o) begin
		main_genericstandalone_crc_errors_status <= (main_genericstandalone_crc_errors_status + 1'd1);
	end
	main_genericstandalone_ps_preamble_error_toggle_o_r <= main_genericstandalone_ps_preamble_error_toggle_o;
	main_genericstandalone_ps_crc_error_toggle_o_r <= main_genericstandalone_ps_crc_error_toggle_o;
	main_genericstandalone_tx_cdc_graycounter0_q_binary <= main_genericstandalone_tx_cdc_graycounter0_q_next_binary;
	main_genericstandalone_tx_cdc_graycounter0_q <= main_genericstandalone_tx_cdc_graycounter0_q_next;
	main_genericstandalone_rx_cdc_graycounter1_q_binary <= main_genericstandalone_rx_cdc_graycounter1_q_next_binary;
	main_genericstandalone_rx_cdc_graycounter1_q <= main_genericstandalone_rx_cdc_graycounter1_q_next;
	if (main_genericstandalone_sram34_counter_reset) begin
		main_genericstandalone_sram33_counter <= 1'd0;
	end else begin
		if (main_genericstandalone_sram35_counter_ce) begin
			main_genericstandalone_sram33_counter <= (main_genericstandalone_sram33_counter + main_genericstandalone_decoded);
		end
	end
	if (main_genericstandalone_slot_ce) begin
		main_genericstandalone_slot <= (main_genericstandalone_slot + 1'd1);
	end
	if (((main_genericstandalone_sram49_we & main_genericstandalone_sram50_writable) & (~main_genericstandalone_sram56_replace))) begin
		main_genericstandalone_sram57_produce <= (main_genericstandalone_sram57_produce + 1'd1);
	end
	if (main_genericstandalone_sram63_do_read) begin
		main_genericstandalone_sram58_consume <= (main_genericstandalone_sram58_consume + 1'd1);
	end
	if (((main_genericstandalone_sram49_we & main_genericstandalone_sram50_writable) & (~main_genericstandalone_sram56_replace))) begin
		if ((~main_genericstandalone_sram63_do_read)) begin
			main_genericstandalone_sram55_level <= (main_genericstandalone_sram55_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_sram63_do_read) begin
			main_genericstandalone_sram55_level <= (main_genericstandalone_sram55_level - 1'd1);
		end
	end
	builder_liteethmacsramwriter_state <= builder_liteethmacsramwriter_next_state;
	if (main_genericstandalone_sram17_status_liteethmac_next_value_ce) begin
		main_genericstandalone_sram17_status <= main_genericstandalone_sram17_status_liteethmac_next_value;
	end
	if (main_genericstandalone_sram153_counter_reset) begin
		main_genericstandalone_sram152_counter <= 1'd0;
	end else begin
		if (main_genericstandalone_sram154_counter_ce) begin
			main_genericstandalone_sram152_counter <= (main_genericstandalone_sram152_counter + 4'd8);
		end
	end
	main_genericstandalone_last_d <= main_genericstandalone_last;
	if (main_genericstandalone_sram109_clear) begin
		main_genericstandalone_sram107_pending <= 1'd0;
	end
	if (main_genericstandalone_sram108_trigger) begin
		main_genericstandalone_sram107_pending <= 1'd1;
	end
	if (((main_genericstandalone_sram129_we & main_genericstandalone_sram130_writable) & (~main_genericstandalone_sram136_replace))) begin
		main_genericstandalone_sram137_produce <= (main_genericstandalone_sram137_produce + 1'd1);
	end
	if (main_genericstandalone_sram143_do_read) begin
		main_genericstandalone_sram138_consume <= (main_genericstandalone_sram138_consume + 1'd1);
	end
	if (((main_genericstandalone_sram129_we & main_genericstandalone_sram130_writable) & (~main_genericstandalone_sram136_replace))) begin
		if ((~main_genericstandalone_sram143_do_read)) begin
			main_genericstandalone_sram135_level <= (main_genericstandalone_sram135_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_sram143_do_read) begin
			main_genericstandalone_sram135_level <= (main_genericstandalone_sram135_level - 1'd1);
		end
	end
	builder_liteethmacsramreader_state <= builder_liteethmacsramreader_next_state;
	main_genericstandalone_sram0_bus_ack <= 1'd0;
	if (((main_genericstandalone_sram0_bus_cyc & main_genericstandalone_sram0_bus_stb) & (~main_genericstandalone_sram0_bus_ack))) begin
		main_genericstandalone_sram0_bus_ack <= 1'd1;
	end
	main_genericstandalone_sram1_bus_ack <= 1'd0;
	if (((main_genericstandalone_sram1_bus_cyc & main_genericstandalone_sram1_bus_stb) & (~main_genericstandalone_sram1_bus_ack))) begin
		main_genericstandalone_sram1_bus_ack <= 1'd1;
	end
	main_genericstandalone_sram2_bus_ack <= 1'd0;
	if (((main_genericstandalone_sram2_bus_cyc & main_genericstandalone_sram2_bus_stb) & (~main_genericstandalone_sram2_bus_ack))) begin
		main_genericstandalone_sram2_bus_ack <= 1'd1;
	end
	main_genericstandalone_sram3_bus_ack <= 1'd0;
	if (((main_genericstandalone_sram3_bus_cyc & main_genericstandalone_sram3_bus_stb) & (~main_genericstandalone_sram3_bus_ack))) begin
		main_genericstandalone_sram3_bus_ack <= 1'd1;
	end
	main_genericstandalone_sram4_bus_ack <= 1'd0;
	if (((main_genericstandalone_sram4_bus_cyc & main_genericstandalone_sram4_bus_stb) & (~main_genericstandalone_sram4_bus_ack))) begin
		main_genericstandalone_sram4_bus_ack <= 1'd1;
	end
	main_genericstandalone_sram5_bus_ack <= 1'd0;
	if (((main_genericstandalone_sram5_bus_cyc & main_genericstandalone_sram5_bus_stb) & (~main_genericstandalone_sram5_bus_ack))) begin
		main_genericstandalone_sram5_bus_ack <= 1'd1;
	end
	main_genericstandalone_sram6_bus_ack <= 1'd0;
	if (((main_genericstandalone_sram6_bus_cyc & main_genericstandalone_sram6_bus_stb) & (~main_genericstandalone_sram6_bus_ack))) begin
		main_genericstandalone_sram6_bus_ack <= 1'd1;
	end
	main_genericstandalone_sram7_bus_ack <= 1'd0;
	if (((main_genericstandalone_sram7_bus_cyc & main_genericstandalone_sram7_bus_stb) & (~main_genericstandalone_sram7_bus_ack))) begin
		main_genericstandalone_sram7_bus_ack <= 1'd1;
	end
	main_genericstandalone_slave_sel_r <= main_genericstandalone_slave_sel;
	case (builder_grant)
		1'd0: begin
			if ((~builder_request[0])) begin
				if (builder_request[1]) begin
					builder_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_request[1])) begin
				if (builder_request[0]) begin
					builder_grant <= 1'd0;
				end
			end
		end
	endcase
	builder_slave_sel_r <= builder_slave_sel;
	main_genericstandalone_mailbox_i1_dat_r <= builder_sync_rhs_self5;
	main_genericstandalone_mailbox_i1_ack <= 1'd0;
	if (((main_genericstandalone_mailbox_i1_cyc & main_genericstandalone_mailbox_i1_stb) & (~main_genericstandalone_mailbox_i1_ack))) begin
		main_genericstandalone_mailbox_i1_ack <= 1'd1;
		if (main_genericstandalone_mailbox_i1_we) begin
			builder_sync_t_t_self0 = main_genericstandalone_mailbox_i1_dat_w;
			case (main_genericstandalone_mailbox_i1_adr[1:0])
				1'd0: begin
					main_genericstandalone_mailbox0 <= builder_sync_t_t_self0;
				end
				1'd1: begin
					main_genericstandalone_mailbox1 <= builder_sync_t_t_self0;
				end
				default: begin
					main_genericstandalone_mailbox2 <= builder_sync_t_t_self0;
				end
			endcase
		end
	end
	main_genericstandalone_mailbox_i2_dat_r <= builder_sync_rhs_self6;
	main_genericstandalone_mailbox_i2_ack <= 1'd0;
	if (((main_genericstandalone_mailbox_i2_cyc & main_genericstandalone_mailbox_i2_stb) & (~main_genericstandalone_mailbox_i2_ack))) begin
		main_genericstandalone_mailbox_i2_ack <= 1'd1;
		if (main_genericstandalone_mailbox_i2_we) begin
			builder_sync_t_t_self1 = main_genericstandalone_mailbox_i2_dat_w;
			case (main_genericstandalone_mailbox_i2_adr[1:0])
				1'd0: begin
					main_genericstandalone_mailbox0 <= builder_sync_t_t_self1;
				end
				1'd1: begin
					main_genericstandalone_mailbox1 <= builder_sync_t_t_self1;
				end
				default: begin
					main_genericstandalone_mailbox2 <= builder_sync_t_t_self1;
				end
			endcase
		end
	end
	if (main_genericstandalone_load) begin
		main_genericstandalone_coarse_ts <= main_genericstandalone_load_value;
	end else begin
		main_genericstandalone_coarse_ts <= (main_genericstandalone_coarse_ts + 1'd1);
	end
	main_genericstandalone_rtio_core_cmd_reset <= main_genericstandalone_rtio_core_reset_re;
	main_genericstandalone_rtio_core_cmd_reset_phy <= main_genericstandalone_rtio_core_reset_phy_re;
	main_genericstandalone_rtio_core_sed_lane_dist_minimum_coarse_timestamp <= (main_genericstandalone_coarse_ts + 4'd12);
	if (main_genericstandalone_rtio_core_async_error_re) begin
		if (main_genericstandalone_rtio_core_async_error_r[0]) begin
			main_genericstandalone_rtio_core_o_collision <= 1'd0;
		end
		if (main_genericstandalone_rtio_core_async_error_r[1]) begin
			main_genericstandalone_rtio_core_o_busy <= 1'd0;
		end
		if (main_genericstandalone_rtio_core_async_error_r[2]) begin
			main_genericstandalone_rtio_core_o_sequence_error <= 1'd0;
		end
	end
	if (main_genericstandalone_rtio_core_o_collision_sync_o) begin
		main_genericstandalone_rtio_core_o_collision <= 1'd1;
		if ((~main_genericstandalone_rtio_core_o_collision)) begin
			main_genericstandalone_rtio_core_collision_channel_status <= main_genericstandalone_rtio_core_o_collision_sync_data_o;
		end
	end
	if (main_genericstandalone_rtio_core_o_busy_sync_o) begin
		main_genericstandalone_rtio_core_o_busy <= 1'd1;
		if ((~main_genericstandalone_rtio_core_o_busy)) begin
			main_genericstandalone_rtio_core_busy_channel_status <= main_genericstandalone_rtio_core_o_busy_sync_data_o;
		end
	end
	if (main_genericstandalone_rtio_core_sed_lane_dist_sequence_error) begin
		main_genericstandalone_rtio_core_o_sequence_error <= 1'd1;
		if ((~main_genericstandalone_rtio_core_o_sequence_error)) begin
			main_genericstandalone_rtio_core_sequence_error_channel_status <= main_genericstandalone_rtio_core_sed_lane_dist_sequence_error_channel;
		end
	end
	main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_o_r <= main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_o;
	if (main_genericstandalone_rtio_core_o_collision_sync_ps_ack_i) begin
		main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_i <= (~main_genericstandalone_rtio_core_o_collision_sync_ps_ack_toggle_i);
	end
	main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_o_r <= main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_o;
	if (main_genericstandalone_rtio_core_o_busy_sync_ps_ack_i) begin
		main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_i <= (~main_genericstandalone_rtio_core_o_busy_sync_ps_ack_toggle_i);
	end
	if (main_genericstandalone_rtio_now_hi_re) begin
		main_genericstandalone_rtio_now_hi_backing <= main_genericstandalone_rtio_now_hi_r;
	end
	if (main_genericstandalone_rtio_now_lo_re) begin
		main_genericstandalone_rtio_now <= {main_genericstandalone_rtio_now_hi_backing, main_genericstandalone_rtio_now_lo_r};
	end
	if (main_genericstandalone_rtio_counter_update_re) begin
		main_genericstandalone_rtio_counter_status <= main_genericstandalone_full_ts;
	end
	case (main_genericstandalone_interface0_csr_bus_adr[4:0])
		1'd0: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_target0_w;
		end
		1'd1: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_rtio_now_hi_w;
		end
		2'd2: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_rtio_now_lo_w;
		end
		2'd3: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data15_w;
		end
		3'd4: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data14_w;
		end
		3'd5: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data13_w;
		end
		3'd6: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data12_w;
		end
		3'd7: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data11_w;
		end
		4'd8: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data10_w;
		end
		4'd9: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data9_w;
		end
		4'd10: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data8_w;
		end
		4'd11: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data7_w;
		end
		4'd12: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data6_w;
		end
		4'd13: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data5_w;
		end
		4'd14: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data4_w;
		end
		4'd15: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data3_w;
		end
		5'd16: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data2_w;
		end
		5'd17: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data1_w;
		end
		5'd18: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_data0_w;
		end
		5'd19: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_o_status_w;
		end
		5'd20: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_i_timeout1_w;
		end
		5'd21: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_i_timeout0_w;
		end
		5'd22: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_i_data_w;
		end
		5'd23: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_i_timestamp1_w;
		end
		5'd24: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_i_timestamp0_w;
		end
		5'd25: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_i_status_w;
		end
		5'd26: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_counter1_w;
		end
		5'd27: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_counter0_w;
		end
		5'd28: begin
			main_genericstandalone_interface0_csr_bus_dat_r <= main_genericstandalone_rtio_counter_update_w;
		end
	endcase
	if (main_genericstandalone_interface0_csr_bus_ack) begin
		main_genericstandalone_interface0_csr_bus_ack <= 1'd0;
	end else begin
		if ((main_genericstandalone_interface0_csr_bus_cyc & main_genericstandalone_interface0_csr_bus_stb)) begin
			main_genericstandalone_interface0_csr_bus_ack <= 1'd1;
		end
	end
	if (main_genericstandalone_target0_re) begin
		main_genericstandalone_rtio_target_storage_full[31:0] <= main_genericstandalone_target0_r;
	end
	main_genericstandalone_rtio_target_re <= main_genericstandalone_target0_re;
	if (main_genericstandalone_rtio_o_data_we) begin
		main_genericstandalone_rtio_o_data_storage_full <= (main_genericstandalone_rtio_o_data_dat_w <<< 1'd0);
	end
	if (main_genericstandalone_o_data15_re) begin
		main_genericstandalone_rtio_o_data_storage_full[511:480] <= main_genericstandalone_o_data15_r;
	end
	if (main_genericstandalone_o_data14_re) begin
		main_genericstandalone_rtio_o_data_storage_full[479:448] <= main_genericstandalone_o_data14_r;
	end
	if (main_genericstandalone_o_data13_re) begin
		main_genericstandalone_rtio_o_data_storage_full[447:416] <= main_genericstandalone_o_data13_r;
	end
	if (main_genericstandalone_o_data12_re) begin
		main_genericstandalone_rtio_o_data_storage_full[415:384] <= main_genericstandalone_o_data12_r;
	end
	if (main_genericstandalone_o_data11_re) begin
		main_genericstandalone_rtio_o_data_storage_full[383:352] <= main_genericstandalone_o_data11_r;
	end
	if (main_genericstandalone_o_data10_re) begin
		main_genericstandalone_rtio_o_data_storage_full[351:320] <= main_genericstandalone_o_data10_r;
	end
	if (main_genericstandalone_o_data9_re) begin
		main_genericstandalone_rtio_o_data_storage_full[319:288] <= main_genericstandalone_o_data9_r;
	end
	if (main_genericstandalone_o_data8_re) begin
		main_genericstandalone_rtio_o_data_storage_full[287:256] <= main_genericstandalone_o_data8_r;
	end
	if (main_genericstandalone_o_data7_re) begin
		main_genericstandalone_rtio_o_data_storage_full[255:224] <= main_genericstandalone_o_data7_r;
	end
	if (main_genericstandalone_o_data6_re) begin
		main_genericstandalone_rtio_o_data_storage_full[223:192] <= main_genericstandalone_o_data6_r;
	end
	if (main_genericstandalone_o_data5_re) begin
		main_genericstandalone_rtio_o_data_storage_full[191:160] <= main_genericstandalone_o_data5_r;
	end
	if (main_genericstandalone_o_data4_re) begin
		main_genericstandalone_rtio_o_data_storage_full[159:128] <= main_genericstandalone_o_data4_r;
	end
	if (main_genericstandalone_o_data3_re) begin
		main_genericstandalone_rtio_o_data_storage_full[127:96] <= main_genericstandalone_o_data3_r;
	end
	if (main_genericstandalone_o_data2_re) begin
		main_genericstandalone_rtio_o_data_storage_full[95:64] <= main_genericstandalone_o_data2_r;
	end
	if (main_genericstandalone_o_data1_re) begin
		main_genericstandalone_rtio_o_data_storage_full[63:32] <= main_genericstandalone_o_data1_r;
	end
	if (main_genericstandalone_o_data0_re) begin
		main_genericstandalone_rtio_o_data_storage_full[31:0] <= main_genericstandalone_o_data0_r;
	end
	main_genericstandalone_rtio_o_data_re <= main_genericstandalone_o_data0_re;
	if (main_genericstandalone_i_timeout1_re) begin
		main_genericstandalone_rtio_i_timeout_storage_full[63:32] <= main_genericstandalone_i_timeout1_r;
	end
	if (main_genericstandalone_i_timeout0_re) begin
		main_genericstandalone_rtio_i_timeout_storage_full[31:0] <= main_genericstandalone_i_timeout0_r;
	end
	main_genericstandalone_rtio_i_timeout_re <= main_genericstandalone_i_timeout0_re;
	case (main_genericstandalone_interface1_csr_bus_adr[3:0])
		1'd0: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_dma_enable_enable_w;
		end
		1'd1: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_base_address1_w;
		end
		2'd2: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_base_address0_w;
		end
		2'd3: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_time_offset1_w;
		end
		3'd4: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_time_offset0_w;
		end
		3'd5: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_dma_cri_master_error_w;
		end
		3'd6: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_error_channel_w;
		end
		3'd7: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_error_timestamp1_w;
		end
		4'd8: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_error_timestamp0_w;
		end
		4'd9: begin
			main_genericstandalone_interface1_csr_bus_dat_r <= main_genericstandalone_error_address_w;
		end
	endcase
	if (main_genericstandalone_interface1_csr_bus_ack) begin
		main_genericstandalone_interface1_csr_bus_ack <= 1'd0;
	end else begin
		if ((main_genericstandalone_interface1_csr_bus_cyc & main_genericstandalone_interface1_csr_bus_stb)) begin
			main_genericstandalone_interface1_csr_bus_ack <= 1'd1;
		end
	end
	if (main_genericstandalone_base_address1_re) begin
		main_genericstandalone_dma_dma_storage_full[32] <= main_genericstandalone_base_address1_r;
	end
	if (main_genericstandalone_base_address0_re) begin
		main_genericstandalone_dma_dma_storage_full[31:0] <= main_genericstandalone_base_address0_r;
	end
	main_genericstandalone_dma_dma_re <= main_genericstandalone_base_address0_re;
	if (main_genericstandalone_time_offset1_re) begin
		main_genericstandalone_dma_time_offset_storage_full[63:32] <= main_genericstandalone_time_offset1_r;
	end
	if (main_genericstandalone_time_offset0_re) begin
		main_genericstandalone_dma_time_offset_storage_full[31:0] <= main_genericstandalone_time_offset0_r;
	end
	main_genericstandalone_dma_time_offset_re <= main_genericstandalone_time_offset0_re;
	main_genericstandalone_cri_con_selected <= main_genericstandalone_cri_con_shared_chan_sel[23:16];
	case (main_genericstandalone_interface2_csr_bus_adr[0])
		1'd0: begin
			main_genericstandalone_interface2_csr_bus_dat_r <= main_genericstandalone_selected0_w;
		end
	endcase
	if (main_genericstandalone_interface2_csr_bus_ack) begin
		main_genericstandalone_interface2_csr_bus_ack <= 1'd0;
	end else begin
		if ((main_genericstandalone_interface2_csr_bus_cyc & main_genericstandalone_interface2_csr_bus_stb)) begin
			main_genericstandalone_interface2_csr_bus_ack <= 1'd1;
		end
	end
	if (main_genericstandalone_selected0_re) begin
		main_genericstandalone_cri_con_storage_full[1:0] <= main_genericstandalone_selected0_r;
	end
	main_genericstandalone_cri_con_re <= main_genericstandalone_selected0_re;
	if (main_genericstandalone_mon_value_update_re) begin
		main_genericstandalone_mon_status <= builder_sync_t_rhs_self3;
	end
	main_genericstandalone_mon_bussynchronizer20_ping_o1 <= main_genericstandalone_mon_bussynchronizer20_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer20_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer20_o <= main_genericstandalone_mon_bussynchronizer20_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer20_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer20_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer20_pong_i) begin
		main_genericstandalone_mon_bussynchronizer20_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer20_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer21_ping_o1 <= main_genericstandalone_mon_bussynchronizer21_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer21_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer21_o <= main_genericstandalone_mon_bussynchronizer21_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer21_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer21_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer21_pong_i) begin
		main_genericstandalone_mon_bussynchronizer21_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer21_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer22_ping_o1 <= main_genericstandalone_mon_bussynchronizer22_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer22_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer22_o <= main_genericstandalone_mon_bussynchronizer22_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer22_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer22_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer22_pong_i) begin
		main_genericstandalone_mon_bussynchronizer22_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer22_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer23_ping_o1 <= main_genericstandalone_mon_bussynchronizer23_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer23_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer23_o <= main_genericstandalone_mon_bussynchronizer23_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer23_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer23_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer23_pong_i) begin
		main_genericstandalone_mon_bussynchronizer23_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer23_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer29_ping_o1 <= main_genericstandalone_mon_bussynchronizer29_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer29_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer29_o <= main_genericstandalone_mon_bussynchronizer29_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer29_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer29_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer29_pong_i) begin
		main_genericstandalone_mon_bussynchronizer29_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer29_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer30_ping_o1 <= main_genericstandalone_mon_bussynchronizer30_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer30_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer30_o <= main_genericstandalone_mon_bussynchronizer30_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer30_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer30_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer30_pong_i) begin
		main_genericstandalone_mon_bussynchronizer30_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer30_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer31_ping_o1 <= main_genericstandalone_mon_bussynchronizer31_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer31_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer31_o <= main_genericstandalone_mon_bussynchronizer31_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer31_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer31_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer31_pong_i) begin
		main_genericstandalone_mon_bussynchronizer31_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer31_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer32_ping_o1 <= main_genericstandalone_mon_bussynchronizer32_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer32_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer32_o <= main_genericstandalone_mon_bussynchronizer32_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer32_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer32_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer32_pong_i) begin
		main_genericstandalone_mon_bussynchronizer32_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer32_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer39_ping_o1 <= main_genericstandalone_mon_bussynchronizer39_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer39_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer39_o <= main_genericstandalone_mon_bussynchronizer39_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer39_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer39_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer39_pong_i) begin
		main_genericstandalone_mon_bussynchronizer39_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer39_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer40_ping_o1 <= main_genericstandalone_mon_bussynchronizer40_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer40_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer40_o <= main_genericstandalone_mon_bussynchronizer40_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer40_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer40_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer40_pong_i) begin
		main_genericstandalone_mon_bussynchronizer40_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer40_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer41_ping_o1 <= main_genericstandalone_mon_bussynchronizer41_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer41_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer41_o <= main_genericstandalone_mon_bussynchronizer41_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer41_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer41_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer41_pong_i) begin
		main_genericstandalone_mon_bussynchronizer41_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer41_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer42_ping_o1 <= main_genericstandalone_mon_bussynchronizer42_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer42_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer42_o <= main_genericstandalone_mon_bussynchronizer42_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer42_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer42_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer42_pong_i) begin
		main_genericstandalone_mon_bussynchronizer42_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer42_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer43_ping_o1 <= main_genericstandalone_mon_bussynchronizer43_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer43_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer43_o <= main_genericstandalone_mon_bussynchronizer43_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer43_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer43_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer43_pong_i) begin
		main_genericstandalone_mon_bussynchronizer43_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer43_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer44_ping_o1 <= main_genericstandalone_mon_bussynchronizer44_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer44_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer44_o <= main_genericstandalone_mon_bussynchronizer44_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer44_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer44_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer44_pong_i) begin
		main_genericstandalone_mon_bussynchronizer44_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer44_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer45_ping_o1 <= main_genericstandalone_mon_bussynchronizer45_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer45_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer45_o <= main_genericstandalone_mon_bussynchronizer45_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer45_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer45_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer45_pong_i) begin
		main_genericstandalone_mon_bussynchronizer45_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer45_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer46_ping_o1 <= main_genericstandalone_mon_bussynchronizer46_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer46_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer46_o <= main_genericstandalone_mon_bussynchronizer46_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer46_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer46_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer46_pong_i) begin
		main_genericstandalone_mon_bussynchronizer46_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer46_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer47_ping_o1 <= main_genericstandalone_mon_bussynchronizer47_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer47_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer47_o <= main_genericstandalone_mon_bussynchronizer47_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer47_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer47_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer47_pong_i) begin
		main_genericstandalone_mon_bussynchronizer47_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer47_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer48_ping_o1 <= main_genericstandalone_mon_bussynchronizer48_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer48_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer48_o <= main_genericstandalone_mon_bussynchronizer48_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer48_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer48_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer48_pong_i) begin
		main_genericstandalone_mon_bussynchronizer48_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer48_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer49_ping_o1 <= main_genericstandalone_mon_bussynchronizer49_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer49_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer49_o <= main_genericstandalone_mon_bussynchronizer49_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer49_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer49_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer49_pong_i) begin
		main_genericstandalone_mon_bussynchronizer49_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer49_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer50_ping_o1 <= main_genericstandalone_mon_bussynchronizer50_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer50_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer50_o <= main_genericstandalone_mon_bussynchronizer50_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer50_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer50_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer50_pong_i) begin
		main_genericstandalone_mon_bussynchronizer50_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer50_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer51_ping_o1 <= main_genericstandalone_mon_bussynchronizer51_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer51_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer51_o <= main_genericstandalone_mon_bussynchronizer51_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer51_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer51_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer51_pong_i) begin
		main_genericstandalone_mon_bussynchronizer51_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer51_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer52_ping_o1 <= main_genericstandalone_mon_bussynchronizer52_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer52_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer52_o <= main_genericstandalone_mon_bussynchronizer52_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer52_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer52_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer52_pong_i) begin
		main_genericstandalone_mon_bussynchronizer52_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer52_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer53_ping_o1 <= main_genericstandalone_mon_bussynchronizer53_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer53_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer53_o <= main_genericstandalone_mon_bussynchronizer53_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer53_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer53_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer53_pong_i) begin
		main_genericstandalone_mon_bussynchronizer53_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer53_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer54_ping_o1 <= main_genericstandalone_mon_bussynchronizer54_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer54_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer54_o <= main_genericstandalone_mon_bussynchronizer54_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer54_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer54_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer54_pong_i) begin
		main_genericstandalone_mon_bussynchronizer54_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer54_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer55_ping_o1 <= main_genericstandalone_mon_bussynchronizer55_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer55_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer55_o <= main_genericstandalone_mon_bussynchronizer55_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer55_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer55_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer55_pong_i) begin
		main_genericstandalone_mon_bussynchronizer55_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer55_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer56_ping_o1 <= main_genericstandalone_mon_bussynchronizer56_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer56_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer56_o <= main_genericstandalone_mon_bussynchronizer56_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer56_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer56_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer56_pong_i) begin
		main_genericstandalone_mon_bussynchronizer56_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer56_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer57_ping_o1 <= main_genericstandalone_mon_bussynchronizer57_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer57_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer57_o <= main_genericstandalone_mon_bussynchronizer57_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer57_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer57_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer57_pong_i) begin
		main_genericstandalone_mon_bussynchronizer57_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer57_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer58_ping_o1 <= main_genericstandalone_mon_bussynchronizer58_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer58_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer58_o <= main_genericstandalone_mon_bussynchronizer58_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer58_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer58_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer58_pong_i) begin
		main_genericstandalone_mon_bussynchronizer58_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer58_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer59_ping_o1 <= main_genericstandalone_mon_bussynchronizer59_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer59_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer59_o <= main_genericstandalone_mon_bussynchronizer59_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer59_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer59_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer59_pong_i) begin
		main_genericstandalone_mon_bussynchronizer59_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer59_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer60_ping_o1 <= main_genericstandalone_mon_bussynchronizer60_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer60_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer60_o <= main_genericstandalone_mon_bussynchronizer60_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer60_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer60_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer60_pong_i) begin
		main_genericstandalone_mon_bussynchronizer60_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer60_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer61_ping_o1 <= main_genericstandalone_mon_bussynchronizer61_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer61_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer61_o <= main_genericstandalone_mon_bussynchronizer61_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer61_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer61_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer61_pong_i) begin
		main_genericstandalone_mon_bussynchronizer61_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer61_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer62_ping_o1 <= main_genericstandalone_mon_bussynchronizer62_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer62_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer62_o <= main_genericstandalone_mon_bussynchronizer62_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer62_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer62_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer62_pong_i) begin
		main_genericstandalone_mon_bussynchronizer62_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer62_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer63_ping_o1 <= main_genericstandalone_mon_bussynchronizer63_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer63_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer63_o <= main_genericstandalone_mon_bussynchronizer63_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer63_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer63_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer63_pong_i) begin
		main_genericstandalone_mon_bussynchronizer63_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer63_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer64_ping_o1 <= main_genericstandalone_mon_bussynchronizer64_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer64_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer64_o <= main_genericstandalone_mon_bussynchronizer64_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer64_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer64_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer64_pong_i) begin
		main_genericstandalone_mon_bussynchronizer64_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer64_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer65_ping_o1 <= main_genericstandalone_mon_bussynchronizer65_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer65_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer65_o <= main_genericstandalone_mon_bussynchronizer65_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer65_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer65_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer65_pong_i) begin
		main_genericstandalone_mon_bussynchronizer65_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer65_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer66_ping_o1 <= main_genericstandalone_mon_bussynchronizer66_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer66_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer66_o <= main_genericstandalone_mon_bussynchronizer66_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer66_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer66_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer66_pong_i) begin
		main_genericstandalone_mon_bussynchronizer66_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer66_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer67_ping_o1 <= main_genericstandalone_mon_bussynchronizer67_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer67_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer67_o <= main_genericstandalone_mon_bussynchronizer67_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer67_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer67_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer67_pong_i) begin
		main_genericstandalone_mon_bussynchronizer67_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer67_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer68_ping_o1 <= main_genericstandalone_mon_bussynchronizer68_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer68_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer68_o <= main_genericstandalone_mon_bussynchronizer68_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer68_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer68_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer68_pong_i) begin
		main_genericstandalone_mon_bussynchronizer68_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer68_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer69_ping_o1 <= main_genericstandalone_mon_bussynchronizer69_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer69_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer69_o <= main_genericstandalone_mon_bussynchronizer69_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer69_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer69_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer69_pong_i) begin
		main_genericstandalone_mon_bussynchronizer69_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer69_pong_toggle_i);
	end
	main_genericstandalone_mon_bussynchronizer70_ping_o1 <= main_genericstandalone_mon_bussynchronizer70_ping_o0;
	if (main_genericstandalone_mon_bussynchronizer70_ping_o1) begin
		main_genericstandalone_mon_bussynchronizer70_o <= main_genericstandalone_mon_bussynchronizer70_obuffer;
	end
	main_genericstandalone_mon_bussynchronizer70_ping_toggle_o_r <= main_genericstandalone_mon_bussynchronizer70_ping_toggle_o;
	if (main_genericstandalone_mon_bussynchronizer70_pong_i) begin
		main_genericstandalone_mon_bussynchronizer70_pong_toggle_i <= (~main_genericstandalone_mon_bussynchronizer70_pong_toggle_i);
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 1'd0)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys0 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 1'd0)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys1 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 1'd0)) & (main_genericstandalone_inj_override_sel_storage == 2'd2))) begin
		main_genericstandalone_inj_o_sys2 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 1'd1)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys3 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 1'd1)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys4 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 1'd1)) & (main_genericstandalone_inj_override_sel_storage == 2'd2))) begin
		main_genericstandalone_inj_o_sys5 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 2'd2)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys6 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 2'd2)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys7 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 2'd2)) & (main_genericstandalone_inj_override_sel_storage == 2'd2))) begin
		main_genericstandalone_inj_o_sys8 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 2'd3)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys9 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 2'd3)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys10 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 2'd3)) & (main_genericstandalone_inj_override_sel_storage == 2'd2))) begin
		main_genericstandalone_inj_o_sys11 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 3'd4)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys12 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 3'd4)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys13 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 3'd5)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys14 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 3'd5)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys15 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 3'd6)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys16 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 3'd6)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys17 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 3'd7)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys18 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 3'd7)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys19 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd8)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys20 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd8)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys21 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd9)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys22 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd9)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys23 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd10)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys24 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd10)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys25 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd11)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys26 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd11)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys27 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd12)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys28 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd12)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys29 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd13)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys30 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd13)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys31 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd14)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys32 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd14)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys33 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd15)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys34 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 4'd15)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys35 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd17)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys36 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd17)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys37 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd18)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys38 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd18)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys39 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd19)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys40 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd19)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys41 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd20)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys42 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd20)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys43 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd21)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys44 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd21)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys45 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd23)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys46 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd23)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys47 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd24)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys48 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd24)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys49 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd25)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys50 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd25)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys51 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd26)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys52 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd26)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys53 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd27)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys54 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd27)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys55 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd30)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys56 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 5'd30)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys57 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd32)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys58 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd32)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys59 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd33)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys60 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd33)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys61 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd34)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys62 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd34)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys63 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd35)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys64 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd35)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys65 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd36)) & (main_genericstandalone_inj_override_sel_storage == 1'd0))) begin
		main_genericstandalone_inj_o_sys66 <= main_genericstandalone_inj_value_r;
	end
	if (((main_genericstandalone_inj_value_re & (main_genericstandalone_inj_chan_sel_storage == 6'd36)) & (main_genericstandalone_inj_override_sel_storage == 1'd1))) begin
		main_genericstandalone_inj_o_sys67 <= main_genericstandalone_inj_value_r;
	end
	main_genericstandalone_rtio_analyzer_enable_r <= main_genericstandalone_rtio_analyzer_enable_storage;
	if ((main_genericstandalone_rtio_analyzer_enable_storage & (~main_genericstandalone_rtio_analyzer_enable_r))) begin
		main_genericstandalone_rtio_analyzer_busy_status <= 1'd1;
	end
	if (((main_genericstandalone_rtio_analyzer_dma_sink_stb & main_genericstandalone_rtio_analyzer_dma_sink_ack) & main_genericstandalone_rtio_analyzer_dma_sink_eop)) begin
		main_genericstandalone_rtio_analyzer_busy_status <= 1'd0;
	end
	main_genericstandalone_rtio_analyzer_message_encoder_read_wait_event_r <= main_genericstandalone_rtio_core_cri_i_status[2];
	main_genericstandalone_rtio_analyzer_message_encoder_just_written <= (main_genericstandalone_rtio_core_cri_cmd == 1'd1);
	main_genericstandalone_rtio_analyzer_message_encoder_enable_r <= main_genericstandalone_rtio_analyzer_enable_storage;
	if (((~main_genericstandalone_rtio_analyzer_enable_storage) & main_genericstandalone_rtio_analyzer_message_encoder_enable_r)) begin
		main_genericstandalone_rtio_analyzer_message_encoder_stopping <= 1'd1;
	end
	if ((~main_genericstandalone_rtio_analyzer_message_encoder_stopping)) begin
		if (main_genericstandalone_rtio_analyzer_message_encoder_exception_stb) begin
			main_genericstandalone_rtio_analyzer_message_encoder_source_payload_data <= {main_genericstandalone_rtio_analyzer_message_encoder_exception_padding1, main_genericstandalone_rtio_analyzer_message_encoder_exception_exception_type, main_genericstandalone_rtio_analyzer_message_encoder_exception_rtio_counter, main_genericstandalone_rtio_analyzer_message_encoder_exception_padding0, main_genericstandalone_rtio_analyzer_message_encoder_exception_channel, main_genericstandalone_rtio_analyzer_message_encoder_exception_message_type};
		end else begin
			main_genericstandalone_rtio_analyzer_message_encoder_source_payload_data <= {main_genericstandalone_rtio_analyzer_message_encoder_input_output_data, main_genericstandalone_rtio_analyzer_message_encoder_input_output_address_padding, main_genericstandalone_rtio_analyzer_message_encoder_input_output_rtio_counter, main_genericstandalone_rtio_analyzer_message_encoder_input_output_timestamp, main_genericstandalone_rtio_analyzer_message_encoder_input_output_channel, main_genericstandalone_rtio_analyzer_message_encoder_input_output_message_type};
		end
		main_genericstandalone_rtio_analyzer_message_encoder_source_eop <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_source_stb <= (main_genericstandalone_rtio_analyzer_enable_storage & (main_genericstandalone_rtio_analyzer_message_encoder_input_output_stb | main_genericstandalone_rtio_analyzer_message_encoder_exception_stb));
		if (main_genericstandalone_rtio_analyzer_message_encoder_overflow_reset_re) begin
			main_genericstandalone_rtio_analyzer_message_encoder_status <= 1'd0;
		end
		if ((main_genericstandalone_rtio_analyzer_message_encoder_source_stb & (~main_genericstandalone_rtio_analyzer_message_encoder_source_ack))) begin
			main_genericstandalone_rtio_analyzer_message_encoder_status <= 1'd1;
		end
	end else begin
		main_genericstandalone_rtio_analyzer_message_encoder_source_payload_data <= {main_genericstandalone_rtio_analyzer_message_encoder_stopped_padding1, main_genericstandalone_rtio_analyzer_message_encoder_stopped_rtio_counter, main_genericstandalone_rtio_analyzer_message_encoder_stopped_padding0, main_genericstandalone_rtio_analyzer_message_encoder_stopped_message_type};
		main_genericstandalone_rtio_analyzer_message_encoder_source_eop <= 1'd1;
		main_genericstandalone_rtio_analyzer_message_encoder_source_stb <= 1'd1;
		if (main_genericstandalone_rtio_analyzer_message_encoder_source_ack) begin
			main_genericstandalone_rtio_analyzer_message_encoder_stopping <= 1'd0;
		end
	end
	if (main_genericstandalone_rtio_analyzer_fifo_transfer_count_rst) begin
		main_genericstandalone_rtio_analyzer_fifo_transfer_count <= 6'd63;
	end else begin
		if (main_genericstandalone_rtio_analyzer_fifo_transfer_count_ce) begin
			main_genericstandalone_rtio_analyzer_fifo_transfer_count <= (main_genericstandalone_rtio_analyzer_fifo_transfer_count - 1'd1);
		end
	end
	main_genericstandalone_rtio_analyzer_fifo_eop_count <= main_genericstandalone_rtio_analyzer_fifo_eop_count_next;
	if ((~main_genericstandalone_rtio_analyzer_fifo_activated)) begin
		main_genericstandalone_rtio_analyzer_fifo_activated <= (main_genericstandalone_rtio_analyzer_fifo_almost_full | (main_genericstandalone_rtio_analyzer_fifo_sink_eop & main_genericstandalone_rtio_analyzer_fifo_do_write));
	end else begin
		if ((main_genericstandalone_rtio_analyzer_fifo_do_read1 & main_genericstandalone_rtio_analyzer_fifo_source_last)) begin
			main_genericstandalone_rtio_analyzer_fifo_activated <= main_genericstandalone_rtio_analyzer_fifo_has_pending_eop;
		end
	end
	if (main_genericstandalone_rtio_analyzer_fifo_syncfifo_re) begin
		main_genericstandalone_rtio_analyzer_fifo_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_rtio_analyzer_fifo_re) begin
			main_genericstandalone_rtio_analyzer_fifo_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_rtio_analyzer_fifo_syncfifo_we & main_genericstandalone_rtio_analyzer_fifo_syncfifo_writable) & (~main_genericstandalone_rtio_analyzer_fifo_replace))) begin
		main_genericstandalone_rtio_analyzer_fifo_produce <= (main_genericstandalone_rtio_analyzer_fifo_produce + 1'd1);
	end
	if (main_genericstandalone_rtio_analyzer_fifo_do_read0) begin
		main_genericstandalone_rtio_analyzer_fifo_consume <= (main_genericstandalone_rtio_analyzer_fifo_consume + 1'd1);
	end
	if (((main_genericstandalone_rtio_analyzer_fifo_syncfifo_we & main_genericstandalone_rtio_analyzer_fifo_syncfifo_writable) & (~main_genericstandalone_rtio_analyzer_fifo_replace))) begin
		if ((~main_genericstandalone_rtio_analyzer_fifo_do_read0)) begin
			main_genericstandalone_rtio_analyzer_fifo_level0 <= (main_genericstandalone_rtio_analyzer_fifo_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_rtio_analyzer_fifo_do_read0) begin
			main_genericstandalone_rtio_analyzer_fifo_level0 <= (main_genericstandalone_rtio_analyzer_fifo_level0 - 1'd1);
		end
	end
	if ((main_genericstandalone_rtio_analyzer_converter_source_stb & main_genericstandalone_rtio_analyzer_converter_source_ack)) begin
		if (main_genericstandalone_rtio_analyzer_converter_last) begin
			main_genericstandalone_rtio_analyzer_converter_mux <= 1'd0;
		end else begin
			main_genericstandalone_rtio_analyzer_converter_mux <= (main_genericstandalone_rtio_analyzer_converter_mux + 1'd1);
		end
	end
	if (main_genericstandalone_rtio_analyzer_dma_reset_re) begin
		main_genericstandalone_interface1_bus_adr <= main_genericstandalone_rtio_analyzer_dma_base_address_storage;
	end
	if (main_genericstandalone_interface1_bus_ack) begin
		if ((main_genericstandalone_interface1_bus_adr == main_genericstandalone_rtio_analyzer_dma_last_address_storage)) begin
			main_genericstandalone_interface1_bus_adr <= main_genericstandalone_rtio_analyzer_dma_base_address_storage;
		end else begin
			main_genericstandalone_interface1_bus_adr <= (main_genericstandalone_interface1_bus_adr + 1'd1);
		end
	end
	if (main_genericstandalone_rtio_analyzer_dma_reset_re) begin
		main_genericstandalone_rtio_analyzer_dma_message_count <= 1'd0;
	end
	if (main_genericstandalone_interface1_bus_ack) begin
		main_genericstandalone_rtio_analyzer_dma_message_count <= (main_genericstandalone_rtio_analyzer_dma_message_count + main_genericstandalone_rtio_analyzer_dma_sink_payload_valid_token_count);
	end
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			if ((~builder_sdram_cpulevel_arbiter_request[0])) begin
				if (builder_sdram_cpulevel_arbiter_request[1]) begin
					builder_sdram_cpulevel_arbiter_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_sdram_cpulevel_arbiter_request[1])) begin
				if (builder_sdram_cpulevel_arbiter_request[0]) begin
					builder_sdram_cpulevel_arbiter_grant <= 1'd0;
				end
			end
		end
	endcase
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			if ((~builder_sdram_native_arbiter_request[0])) begin
				if (builder_sdram_native_arbiter_request[1]) begin
					builder_sdram_native_arbiter_grant <= 1'd1;
				end else begin
					if (builder_sdram_native_arbiter_request[2]) begin
						builder_sdram_native_arbiter_grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~builder_sdram_native_arbiter_request[1])) begin
				if (builder_sdram_native_arbiter_request[2]) begin
					builder_sdram_native_arbiter_grant <= 2'd2;
				end else begin
					if (builder_sdram_native_arbiter_request[0]) begin
						builder_sdram_native_arbiter_grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~builder_sdram_native_arbiter_request[2])) begin
				if (builder_sdram_native_arbiter_request[0]) begin
					builder_sdram_native_arbiter_grant <= 1'd0;
				end else begin
					if (builder_sdram_native_arbiter_request[1]) begin
						builder_sdram_native_arbiter_grant <= 1'd1;
					end
				end
			end
		end
	endcase
	case (builder_genericstandalone_grant)
		1'd0: begin
			if ((~builder_genericstandalone_request[0])) begin
				if (builder_genericstandalone_request[1]) begin
					builder_genericstandalone_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_genericstandalone_request[1])) begin
				if (builder_genericstandalone_request[0]) begin
					builder_genericstandalone_grant <= 1'd0;
				end
			end
		end
	endcase
	builder_genericstandalone_slave_sel_r <= builder_genericstandalone_slave_sel;
	builder_genericstandalone_interface0_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank0_sel) begin
		case (builder_genericstandalone_interface0_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface0_bank_bus_dat_r <= builder_genericstandalone_csrbank0_switch_done_w;
			end
			1'd1: begin
				builder_genericstandalone_interface0_bank_bus_dat_r <= builder_genericstandalone_csrbank0_clock_sel0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank0_clock_sel0_re) begin
		main_genericstandalone_rtiosyscrg_storage_full <= builder_genericstandalone_csrbank0_clock_sel0_r;
	end
	main_genericstandalone_rtiosyscrg_re <= builder_genericstandalone_csrbank0_clock_sel0_re;
	builder_genericstandalone_interface1_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank1_sel) begin
		case (builder_genericstandalone_interface1_bank_bus_adr[1:0])
			1'd0: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_dly_sel0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_w;
			end
			2'd2: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_w;
			end
			2'd3: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank1_dly_sel0_re) begin
		main_genericstandalone_genericstandalone_ddrphy_storage_full[1:0] <= builder_genericstandalone_csrbank1_dly_sel0_r;
	end
	main_genericstandalone_genericstandalone_ddrphy_re <= builder_genericstandalone_csrbank1_dly_sel0_re;
	builder_genericstandalone_interface2_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank2_sel) begin
		case (builder_genericstandalone_interface2_bank_bus_adr[5:0])
			1'd0: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_control0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_command0_w;
			end
			2'd2: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_address1_w;
			end
			3'd4: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_address0_w;
			end
			3'd5: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_baddress0_w;
			end
			3'd6: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_wrdata3_w;
			end
			3'd7: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_wrdata2_w;
			end
			4'd8: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_wrdata1_w;
			end
			4'd9: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_wrdata0_w;
			end
			4'd10: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_rddata3_w;
			end
			4'd11: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_rddata2_w;
			end
			4'd12: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_rddata1_w;
			end
			4'd13: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi0_rddata0_w;
			end
			4'd14: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_command0_w;
			end
			4'd15: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_w;
			end
			5'd16: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_address1_w;
			end
			5'd17: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_address0_w;
			end
			5'd18: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_baddress0_w;
			end
			5'd19: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_wrdata3_w;
			end
			5'd20: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_wrdata2_w;
			end
			5'd21: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_wrdata1_w;
			end
			5'd22: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_wrdata0_w;
			end
			5'd23: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_rddata3_w;
			end
			5'd24: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_rddata2_w;
			end
			5'd25: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_rddata1_w;
			end
			5'd26: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi1_rddata0_w;
			end
			5'd27: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_command0_w;
			end
			5'd28: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_w;
			end
			5'd29: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_address1_w;
			end
			5'd30: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_address0_w;
			end
			5'd31: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_baddress0_w;
			end
			6'd32: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_wrdata3_w;
			end
			6'd33: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_wrdata2_w;
			end
			6'd34: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_wrdata1_w;
			end
			6'd35: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_wrdata0_w;
			end
			6'd36: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_rddata3_w;
			end
			6'd37: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_rddata2_w;
			end
			6'd38: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_rddata1_w;
			end
			6'd39: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi2_rddata0_w;
			end
			6'd40: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_command0_w;
			end
			6'd41: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_w;
			end
			6'd42: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_address1_w;
			end
			6'd43: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_address0_w;
			end
			6'd44: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_baddress0_w;
			end
			6'd45: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_wrdata3_w;
			end
			6'd46: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_wrdata2_w;
			end
			6'd47: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_wrdata1_w;
			end
			6'd48: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_wrdata0_w;
			end
			6'd49: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_rddata3_w;
			end
			6'd50: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_rddata2_w;
			end
			6'd51: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_rddata1_w;
			end
			6'd52: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_pi3_rddata0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank2_control0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_storage_full[3:0] <= builder_genericstandalone_csrbank2_control0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_re <= builder_genericstandalone_csrbank2_control0_re;
	if (builder_genericstandalone_csrbank2_pi0_command0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full[5:0] <= builder_genericstandalone_csrbank2_pi0_command0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_re <= builder_genericstandalone_csrbank2_pi0_command0_re;
	if (builder_genericstandalone_csrbank2_pi0_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[14:8] <= builder_genericstandalone_csrbank2_pi0_address1_r;
	end
	if (builder_genericstandalone_csrbank2_pi0_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[7:0] <= builder_genericstandalone_csrbank2_pi0_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_re <= builder_genericstandalone_csrbank2_pi0_address0_re;
	if (builder_genericstandalone_csrbank2_pi0_baddress0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full[2:0] <= builder_genericstandalone_csrbank2_pi0_baddress0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_re <= builder_genericstandalone_csrbank2_pi0_baddress0_re;
	if (builder_genericstandalone_csrbank2_pi0_wrdata3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[31:24] <= builder_genericstandalone_csrbank2_pi0_wrdata3_r;
	end
	if (builder_genericstandalone_csrbank2_pi0_wrdata2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[23:16] <= builder_genericstandalone_csrbank2_pi0_wrdata2_r;
	end
	if (builder_genericstandalone_csrbank2_pi0_wrdata1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[15:8] <= builder_genericstandalone_csrbank2_pi0_wrdata1_r;
	end
	if (builder_genericstandalone_csrbank2_pi0_wrdata0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[7:0] <= builder_genericstandalone_csrbank2_pi0_wrdata0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_re <= builder_genericstandalone_csrbank2_pi0_wrdata0_re;
	if (builder_genericstandalone_csrbank2_pi1_command0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full[5:0] <= builder_genericstandalone_csrbank2_pi1_command0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_re <= builder_genericstandalone_csrbank2_pi1_command0_re;
	if (builder_genericstandalone_csrbank2_pi1_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[14:8] <= builder_genericstandalone_csrbank2_pi1_address1_r;
	end
	if (builder_genericstandalone_csrbank2_pi1_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[7:0] <= builder_genericstandalone_csrbank2_pi1_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_re <= builder_genericstandalone_csrbank2_pi1_address0_re;
	if (builder_genericstandalone_csrbank2_pi1_baddress0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full[2:0] <= builder_genericstandalone_csrbank2_pi1_baddress0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_re <= builder_genericstandalone_csrbank2_pi1_baddress0_re;
	if (builder_genericstandalone_csrbank2_pi1_wrdata3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[31:24] <= builder_genericstandalone_csrbank2_pi1_wrdata3_r;
	end
	if (builder_genericstandalone_csrbank2_pi1_wrdata2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[23:16] <= builder_genericstandalone_csrbank2_pi1_wrdata2_r;
	end
	if (builder_genericstandalone_csrbank2_pi1_wrdata1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[15:8] <= builder_genericstandalone_csrbank2_pi1_wrdata1_r;
	end
	if (builder_genericstandalone_csrbank2_pi1_wrdata0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[7:0] <= builder_genericstandalone_csrbank2_pi1_wrdata0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_re <= builder_genericstandalone_csrbank2_pi1_wrdata0_re;
	if (builder_genericstandalone_csrbank2_pi2_command0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full[5:0] <= builder_genericstandalone_csrbank2_pi2_command0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_re <= builder_genericstandalone_csrbank2_pi2_command0_re;
	if (builder_genericstandalone_csrbank2_pi2_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[14:8] <= builder_genericstandalone_csrbank2_pi2_address1_r;
	end
	if (builder_genericstandalone_csrbank2_pi2_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[7:0] <= builder_genericstandalone_csrbank2_pi2_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_re <= builder_genericstandalone_csrbank2_pi2_address0_re;
	if (builder_genericstandalone_csrbank2_pi2_baddress0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full[2:0] <= builder_genericstandalone_csrbank2_pi2_baddress0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_re <= builder_genericstandalone_csrbank2_pi2_baddress0_re;
	if (builder_genericstandalone_csrbank2_pi2_wrdata3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[31:24] <= builder_genericstandalone_csrbank2_pi2_wrdata3_r;
	end
	if (builder_genericstandalone_csrbank2_pi2_wrdata2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[23:16] <= builder_genericstandalone_csrbank2_pi2_wrdata2_r;
	end
	if (builder_genericstandalone_csrbank2_pi2_wrdata1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[15:8] <= builder_genericstandalone_csrbank2_pi2_wrdata1_r;
	end
	if (builder_genericstandalone_csrbank2_pi2_wrdata0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[7:0] <= builder_genericstandalone_csrbank2_pi2_wrdata0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_re <= builder_genericstandalone_csrbank2_pi2_wrdata0_re;
	if (builder_genericstandalone_csrbank2_pi3_command0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full[5:0] <= builder_genericstandalone_csrbank2_pi3_command0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_re <= builder_genericstandalone_csrbank2_pi3_command0_re;
	if (builder_genericstandalone_csrbank2_pi3_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[14:8] <= builder_genericstandalone_csrbank2_pi3_address1_r;
	end
	if (builder_genericstandalone_csrbank2_pi3_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[7:0] <= builder_genericstandalone_csrbank2_pi3_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_re <= builder_genericstandalone_csrbank2_pi3_address0_re;
	if (builder_genericstandalone_csrbank2_pi3_baddress0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full[2:0] <= builder_genericstandalone_csrbank2_pi3_baddress0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_re <= builder_genericstandalone_csrbank2_pi3_baddress0_re;
	if (builder_genericstandalone_csrbank2_pi3_wrdata3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[31:24] <= builder_genericstandalone_csrbank2_pi3_wrdata3_r;
	end
	if (builder_genericstandalone_csrbank2_pi3_wrdata2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[23:16] <= builder_genericstandalone_csrbank2_pi3_wrdata2_r;
	end
	if (builder_genericstandalone_csrbank2_pi3_wrdata1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[15:8] <= builder_genericstandalone_csrbank2_pi3_wrdata1_r;
	end
	if (builder_genericstandalone_csrbank2_pi3_wrdata0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[7:0] <= builder_genericstandalone_csrbank2_pi3_wrdata0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_re <= builder_genericstandalone_csrbank2_pi3_wrdata0_re;
	builder_genericstandalone_interface3_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank3_sel) begin
		case (builder_genericstandalone_interface3_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface3_bank_bus_dat_r <= builder_genericstandalone_csrbank3_out0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank3_out0_re) begin
		main_genericstandalone_error_led_storage_full <= builder_genericstandalone_csrbank3_out0_r;
	end
	main_genericstandalone_error_led_re <= builder_genericstandalone_csrbank3_out0_re;
	builder_genericstandalone_interface4_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank4_sel) begin
		case (builder_genericstandalone_interface4_bank_bus_adr[4:0])
			1'd0: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_writer_slot_w;
			end
			1'd1: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_writer_length1_w;
			end
			2'd2: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_writer_length0_w;
			end
			2'd3: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_writer_errors3_w;
			end
			3'd4: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_writer_errors2_w;
			end
			3'd5: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_writer_errors1_w;
			end
			3'd6: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_writer_errors0_w;
			end
			3'd7: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= main_genericstandalone_sram25_status_w;
			end
			4'd8: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= main_genericstandalone_sram28_pending_w;
			end
			4'd9: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_writer_ev_enable0_w;
			end
			4'd10: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= main_genericstandalone_start_w;
			end
			4'd11: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_reader_ready_w;
			end
			4'd12: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_reader_slot0_w;
			end
			4'd13: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_reader_length1_w;
			end
			4'd14: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_reader_length0_w;
			end
			4'd15: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= main_genericstandalone_sram112_status_w;
			end
			5'd16: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= main_genericstandalone_sram115_pending_w;
			end
			5'd17: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_sram_reader_ev_enable0_w;
			end
			5'd18: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_preamble_errors3_w;
			end
			5'd19: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_preamble_errors2_w;
			end
			5'd20: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_preamble_errors1_w;
			end
			5'd21: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_preamble_errors0_w;
			end
			5'd22: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_crc_errors3_w;
			end
			5'd23: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_crc_errors2_w;
			end
			5'd24: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_crc_errors1_w;
			end
			5'd25: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_crc_errors0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank4_sram_writer_ev_enable0_re) begin
		main_genericstandalone_sram29_storage_full <= builder_genericstandalone_csrbank4_sram_writer_ev_enable0_r;
	end
	main_genericstandalone_sram31_re <= builder_genericstandalone_csrbank4_sram_writer_ev_enable0_re;
	if (builder_genericstandalone_csrbank4_sram_reader_slot0_re) begin
		main_genericstandalone_sram99_storage_full[1:0] <= builder_genericstandalone_csrbank4_sram_reader_slot0_r;
	end
	main_genericstandalone_sram101_re <= builder_genericstandalone_csrbank4_sram_reader_slot0_re;
	if (builder_genericstandalone_csrbank4_sram_reader_length1_re) begin
		main_genericstandalone_sram102_storage_full[10:8] <= builder_genericstandalone_csrbank4_sram_reader_length1_r;
	end
	if (builder_genericstandalone_csrbank4_sram_reader_length0_re) begin
		main_genericstandalone_sram102_storage_full[7:0] <= builder_genericstandalone_csrbank4_sram_reader_length0_r;
	end
	main_genericstandalone_sram104_re <= builder_genericstandalone_csrbank4_sram_reader_length0_re;
	if (builder_genericstandalone_csrbank4_sram_reader_ev_enable0_re) begin
		main_genericstandalone_sram116_storage_full <= builder_genericstandalone_csrbank4_sram_reader_ev_enable0_r;
	end
	main_genericstandalone_sram118_re <= builder_genericstandalone_csrbank4_sram_reader_ev_enable0_re;
	builder_genericstandalone_interface5_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank5_sel) begin
		case (builder_genericstandalone_interface5_bank_bus_adr[1:0])
			1'd0: begin
				builder_genericstandalone_interface5_bank_bus_dat_r <= builder_genericstandalone_csrbank5_in_w;
			end
			1'd1: begin
				builder_genericstandalone_interface5_bank_bus_dat_r <= builder_genericstandalone_csrbank5_out0_w;
			end
			2'd2: begin
				builder_genericstandalone_interface5_bank_bus_dat_r <= builder_genericstandalone_csrbank5_oe0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank5_out0_re) begin
		main_genericstandalone_i2c_out_storage_full[1:0] <= builder_genericstandalone_csrbank5_out0_r;
	end
	main_genericstandalone_i2c_out_re <= builder_genericstandalone_csrbank5_out0_re;
	if (builder_genericstandalone_csrbank5_oe0_re) begin
		main_genericstandalone_i2c_oe_storage_full[1:0] <= builder_genericstandalone_csrbank5_oe0_r;
	end
	main_genericstandalone_i2c_oe_re <= builder_genericstandalone_csrbank5_oe0_re;
	builder_genericstandalone_interface6_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank6_sel) begin
		case (builder_genericstandalone_interface6_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface6_bank_bus_dat_r <= main_genericstandalone_genericstandalone_icap_iprog_w;
			end
		endcase
	end
	builder_genericstandalone_interface7_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank7_sel) begin
		case (builder_genericstandalone_interface7_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_address0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_data_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank7_address0_re) begin
		main_genericstandalone_add_identifier_storage_full[7:0] <= builder_genericstandalone_csrbank7_address0_r;
	end
	main_genericstandalone_add_identifier_re <= builder_genericstandalone_csrbank7_address0_re;
	builder_genericstandalone_interface8_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank8_sel) begin
		case (builder_genericstandalone_interface8_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= builder_genericstandalone_csrbank8_reset0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank8_reset0_re) begin
		main_genericstandalone_kernel_cpu_storage_full <= builder_genericstandalone_csrbank8_reset0_r;
	end
	main_genericstandalone_kernel_cpu_re <= builder_genericstandalone_csrbank8_reset0_re;
	builder_genericstandalone_interface9_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank9_sel) begin
		case (builder_genericstandalone_interface9_bank_bus_adr[4:0])
			1'd0: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_enable0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_busy_w;
			end
			2'd2: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_message_encoder_overflow_w;
			end
			2'd3: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= main_genericstandalone_rtio_analyzer_message_encoder_overflow_reset_w;
			end
			3'd4: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= main_genericstandalone_rtio_analyzer_dma_reset_w;
			end
			3'd5: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_base_address4_w;
			end
			3'd6: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_base_address3_w;
			end
			3'd7: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_base_address2_w;
			end
			4'd8: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_base_address1_w;
			end
			4'd9: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_base_address0_w;
			end
			4'd10: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_last_address4_w;
			end
			4'd11: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_last_address3_w;
			end
			4'd12: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_last_address2_w;
			end
			4'd13: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_last_address1_w;
			end
			4'd14: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_last_address0_w;
			end
			4'd15: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_byte_count7_w;
			end
			5'd16: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_byte_count6_w;
			end
			5'd17: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_byte_count5_w;
			end
			5'd18: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_byte_count4_w;
			end
			5'd19: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_byte_count3_w;
			end
			5'd20: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_byte_count2_w;
			end
			5'd21: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_byte_count1_w;
			end
			5'd22: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_dma_byte_count0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank9_enable0_re) begin
		main_genericstandalone_rtio_analyzer_enable_storage_full <= builder_genericstandalone_csrbank9_enable0_r;
	end
	main_genericstandalone_rtio_analyzer_enable_re <= builder_genericstandalone_csrbank9_enable0_re;
	if (builder_genericstandalone_csrbank9_dma_base_address4_re) begin
		main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[32] <= builder_genericstandalone_csrbank9_dma_base_address4_r;
	end
	if (builder_genericstandalone_csrbank9_dma_base_address3_re) begin
		main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[31:24] <= builder_genericstandalone_csrbank9_dma_base_address3_r;
	end
	if (builder_genericstandalone_csrbank9_dma_base_address2_re) begin
		main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[23:16] <= builder_genericstandalone_csrbank9_dma_base_address2_r;
	end
	if (builder_genericstandalone_csrbank9_dma_base_address1_re) begin
		main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[15:8] <= builder_genericstandalone_csrbank9_dma_base_address1_r;
	end
	if (builder_genericstandalone_csrbank9_dma_base_address0_re) begin
		main_genericstandalone_rtio_analyzer_dma_base_address_storage_full[7:0] <= builder_genericstandalone_csrbank9_dma_base_address0_r;
	end
	main_genericstandalone_rtio_analyzer_dma_base_address_re <= builder_genericstandalone_csrbank9_dma_base_address0_re;
	if (builder_genericstandalone_csrbank9_dma_last_address4_re) begin
		main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[32] <= builder_genericstandalone_csrbank9_dma_last_address4_r;
	end
	if (builder_genericstandalone_csrbank9_dma_last_address3_re) begin
		main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[31:24] <= builder_genericstandalone_csrbank9_dma_last_address3_r;
	end
	if (builder_genericstandalone_csrbank9_dma_last_address2_re) begin
		main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[23:16] <= builder_genericstandalone_csrbank9_dma_last_address2_r;
	end
	if (builder_genericstandalone_csrbank9_dma_last_address1_re) begin
		main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[15:8] <= builder_genericstandalone_csrbank9_dma_last_address1_r;
	end
	if (builder_genericstandalone_csrbank9_dma_last_address0_re) begin
		main_genericstandalone_rtio_analyzer_dma_last_address_storage_full[7:0] <= builder_genericstandalone_csrbank9_dma_last_address0_r;
	end
	main_genericstandalone_rtio_analyzer_dma_last_address_re <= builder_genericstandalone_csrbank9_dma_last_address0_re;
	builder_genericstandalone_interface10_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank10_sel) begin
		case (builder_genericstandalone_interface10_bank_bus_adr[3:0])
			1'd0: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= main_genericstandalone_rtio_core_reset_w;
			end
			1'd1: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= main_genericstandalone_rtio_core_reset_phy_w;
			end
			2'd2: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_sed_spread_enable0_w;
			end
			2'd3: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= main_genericstandalone_rtio_core_async_error_w;
			end
			3'd4: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_collision_channel1_w;
			end
			3'd5: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_collision_channel0_w;
			end
			3'd6: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_busy_channel1_w;
			end
			3'd7: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_busy_channel0_w;
			end
			4'd8: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_sequence_error_channel1_w;
			end
			4'd9: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_sequence_error_channel0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank10_sed_spread_enable0_re) begin
		main_genericstandalone_rtio_core_storage_full <= builder_genericstandalone_csrbank10_sed_spread_enable0_r;
	end
	main_genericstandalone_rtio_core_re <= builder_genericstandalone_csrbank10_sed_spread_enable0_re;
	builder_genericstandalone_interface11_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank11_sel) begin
		case (builder_genericstandalone_interface11_bank_bus_adr[3:0])
			1'd0: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_mon_chan_sel0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_mon_probe_sel0_w;
			end
			2'd2: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= main_genericstandalone_mon_value_update_w;
			end
			2'd3: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_mon_value3_w;
			end
			3'd4: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_mon_value2_w;
			end
			3'd5: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_mon_value1_w;
			end
			3'd6: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_mon_value0_w;
			end
			3'd7: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_inj_chan_sel0_w;
			end
			4'd8: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_inj_override_sel0_w;
			end
			4'd9: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= main_genericstandalone_inj_value_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank11_mon_chan_sel0_re) begin
		main_genericstandalone_mon_chan_sel_storage_full[5:0] <= builder_genericstandalone_csrbank11_mon_chan_sel0_r;
	end
	main_genericstandalone_mon_chan_sel_re <= builder_genericstandalone_csrbank11_mon_chan_sel0_re;
	if (builder_genericstandalone_csrbank11_mon_probe_sel0_re) begin
		main_genericstandalone_mon_probe_sel_storage_full[4:0] <= builder_genericstandalone_csrbank11_mon_probe_sel0_r;
	end
	main_genericstandalone_mon_probe_sel_re <= builder_genericstandalone_csrbank11_mon_probe_sel0_re;
	if (builder_genericstandalone_csrbank11_inj_chan_sel0_re) begin
		main_genericstandalone_inj_chan_sel_storage_full[5:0] <= builder_genericstandalone_csrbank11_inj_chan_sel0_r;
	end
	main_genericstandalone_inj_chan_sel_re <= builder_genericstandalone_csrbank11_inj_chan_sel0_re;
	if (builder_genericstandalone_csrbank11_inj_override_sel0_re) begin
		main_genericstandalone_inj_override_sel_storage_full[1:0] <= builder_genericstandalone_csrbank11_inj_override_sel0_r;
	end
	main_genericstandalone_inj_override_sel_re <= builder_genericstandalone_csrbank11_inj_override_sel0_re;
	builder_genericstandalone_interface12_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank12_sel) begin
		case (builder_genericstandalone_interface12_bank_bus_adr[1:0])
			1'd0: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_bitbang0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_miso_w;
			end
			2'd2: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_bitbang_en0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank12_bitbang0_re) begin
		main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full[3:0] <= builder_genericstandalone_csrbank12_bitbang0_r;
	end
	main_genericstandalone_genericstandalone_spiflash_bitbang_re <= builder_genericstandalone_csrbank12_bitbang0_re;
	if (builder_genericstandalone_csrbank12_bitbang_en0_re) begin
		main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full <= builder_genericstandalone_csrbank12_bitbang_en0_r;
	end
	main_genericstandalone_genericstandalone_spiflash_bitbang_en_re <= builder_genericstandalone_csrbank12_bitbang_en0_re;
	builder_genericstandalone_interface13_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank13_sel) begin
		case (builder_genericstandalone_interface13_bank_bus_adr[4:0])
			1'd0: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_load7_w;
			end
			1'd1: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_load6_w;
			end
			2'd2: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_load5_w;
			end
			2'd3: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_load4_w;
			end
			3'd4: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_load3_w;
			end
			3'd5: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_load2_w;
			end
			3'd6: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_load1_w;
			end
			3'd7: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_load0_w;
			end
			4'd8: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_reload7_w;
			end
			4'd9: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_reload6_w;
			end
			4'd10: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_reload5_w;
			end
			4'd11: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_reload4_w;
			end
			4'd12: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_reload3_w;
			end
			4'd13: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_reload2_w;
			end
			4'd14: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_reload1_w;
			end
			4'd15: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_reload0_w;
			end
			5'd16: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_en0_w;
			end
			5'd17: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_w;
			end
			5'd18: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_value7_w;
			end
			5'd19: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_value6_w;
			end
			5'd20: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_value5_w;
			end
			5'd21: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_value4_w;
			end
			5'd22: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_value3_w;
			end
			5'd23: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_value2_w;
			end
			5'd24: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_value1_w;
			end
			5'd25: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_value0_w;
			end
			5'd26: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_w;
			end
			5'd27: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_w;
			end
			5'd28: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_ev_enable0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank13_load7_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[63:56] <= builder_genericstandalone_csrbank13_load7_r;
	end
	if (builder_genericstandalone_csrbank13_load6_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[55:48] <= builder_genericstandalone_csrbank13_load6_r;
	end
	if (builder_genericstandalone_csrbank13_load5_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[47:40] <= builder_genericstandalone_csrbank13_load5_r;
	end
	if (builder_genericstandalone_csrbank13_load4_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[39:32] <= builder_genericstandalone_csrbank13_load4_r;
	end
	if (builder_genericstandalone_csrbank13_load3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[31:24] <= builder_genericstandalone_csrbank13_load3_r;
	end
	if (builder_genericstandalone_csrbank13_load2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[23:16] <= builder_genericstandalone_csrbank13_load2_r;
	end
	if (builder_genericstandalone_csrbank13_load1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[15:8] <= builder_genericstandalone_csrbank13_load1_r;
	end
	if (builder_genericstandalone_csrbank13_load0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[7:0] <= builder_genericstandalone_csrbank13_load0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_load_re <= builder_genericstandalone_csrbank13_load0_re;
	if (builder_genericstandalone_csrbank13_reload7_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[63:56] <= builder_genericstandalone_csrbank13_reload7_r;
	end
	if (builder_genericstandalone_csrbank13_reload6_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[55:48] <= builder_genericstandalone_csrbank13_reload6_r;
	end
	if (builder_genericstandalone_csrbank13_reload5_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[47:40] <= builder_genericstandalone_csrbank13_reload5_r;
	end
	if (builder_genericstandalone_csrbank13_reload4_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[39:32] <= builder_genericstandalone_csrbank13_reload4_r;
	end
	if (builder_genericstandalone_csrbank13_reload3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[31:24] <= builder_genericstandalone_csrbank13_reload3_r;
	end
	if (builder_genericstandalone_csrbank13_reload2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[23:16] <= builder_genericstandalone_csrbank13_reload2_r;
	end
	if (builder_genericstandalone_csrbank13_reload1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[15:8] <= builder_genericstandalone_csrbank13_reload1_r;
	end
	if (builder_genericstandalone_csrbank13_reload0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[7:0] <= builder_genericstandalone_csrbank13_reload0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_re <= builder_genericstandalone_csrbank13_reload0_re;
	if (builder_genericstandalone_csrbank13_en0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full <= builder_genericstandalone_csrbank13_en0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_en_re <= builder_genericstandalone_csrbank13_en0_re;
	if (builder_genericstandalone_csrbank13_ev_enable0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full <= builder_genericstandalone_csrbank13_ev_enable0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_re <= builder_genericstandalone_csrbank13_ev_enable0_re;
	builder_genericstandalone_interface14_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank14_sel) begin
		case (builder_genericstandalone_interface14_bank_bus_adr[2:0])
			1'd0: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_w;
			end
			1'd1: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= builder_genericstandalone_csrbank14_txfull_w;
			end
			2'd2: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= builder_genericstandalone_csrbank14_rxempty_w;
			end
			2'd3: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_uart_status_w;
			end
			3'd4: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w;
			end
			3'd5: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= builder_genericstandalone_csrbank14_ev_enable0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank14_ev_enable0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full[1:0] <= builder_genericstandalone_csrbank14_ev_enable0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_re <= builder_genericstandalone_csrbank14_ev_enable0_re;
	builder_genericstandalone_interface15_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank15_sel) begin
		case (builder_genericstandalone_interface15_bank_bus_adr[1:0])
			1'd0: begin
				builder_genericstandalone_interface15_bank_bus_dat_r <= builder_genericstandalone_csrbank15_tuning_word3_w;
			end
			1'd1: begin
				builder_genericstandalone_interface15_bank_bus_dat_r <= builder_genericstandalone_csrbank15_tuning_word2_w;
			end
			2'd2: begin
				builder_genericstandalone_interface15_bank_bus_dat_r <= builder_genericstandalone_csrbank15_tuning_word1_w;
			end
			2'd3: begin
				builder_genericstandalone_interface15_bank_bus_dat_r <= builder_genericstandalone_csrbank15_tuning_word0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank15_tuning_word3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[31:24] <= builder_genericstandalone_csrbank15_tuning_word3_r;
	end
	if (builder_genericstandalone_csrbank15_tuning_word2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[23:16] <= builder_genericstandalone_csrbank15_tuning_word2_r;
	end
	if (builder_genericstandalone_csrbank15_tuning_word1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[15:8] <= builder_genericstandalone_csrbank15_tuning_word1_r;
	end
	if (builder_genericstandalone_csrbank15_tuning_word0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[7:0] <= builder_genericstandalone_csrbank15_tuning_word0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_phy_re <= builder_genericstandalone_csrbank15_tuning_word0_re;
	builder_genericstandalone_interface16_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank16_sel) begin
		case (builder_genericstandalone_interface16_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface16_bank_bus_dat_r <= builder_genericstandalone_csrbank16_status_w;
			end
		endcase
	end
	if (sys_rst) begin
		main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_interface_adr <= 14'd0;
		main_genericstandalone_genericstandalone_genericstandalone_interface_we <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w <= 8'd0;
		main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_r <= 64'd0;
		main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_trigger <= 2'd0;
		serial_tx <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full <= 32'd3958241;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg <= 8'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_payload_data <= 8'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_r <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg <= 8'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_old_trigger <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_old_trigger <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full <= 2'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level <= 5'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level <= 5'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full <= 64'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full <= 64'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_en_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status <= 64'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_old_trigger <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_value <= 64'd0;
		main_genericstandalone_genericstandalone_ddrphy_storage_full <= 2'd0;
		main_genericstandalone_genericstandalone_ddrphy_re <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_valid <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_valid <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_valid <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_valid <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_oe_dqs <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_oe_dq <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en0 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en1 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en2 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en3 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_storage_full <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full <= 6'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full <= 3'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full <= 6'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full <= 3'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full <= 6'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full <= 3'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full <= 6'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full <= 3'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_mask <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_mask <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_mask <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_mask <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_count <= 3'd4;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_pending_refresh <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refi_cycles <= 10'd977;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_sdram_col <= 10'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_rdvalid_r <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_dat_w0 <= 128'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_sel0 <= 16'd0;
		main_genericstandalone_genericstandalone_genericstandalone_cache <= 2'd0;
		main_genericstandalone_genericstandalone_genericstandalone_cache_adr_offset_r <= 3'd0;
		main_genericstandalone_genericstandalone_spiflash_bus_ack <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full <= 4'd0;
		main_genericstandalone_genericstandalone_spiflash_bitbang_re <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_bitbang_en_re <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_spiflash_clk <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_dq_oe <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_sr <= 64'd0;
		main_genericstandalone_genericstandalone_spiflash_i1 <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_dqi <= 2'd0;
		main_genericstandalone_genericstandalone_spiflash_trigger <= 7'd0;
		main_genericstandalone_tx_mmcm_reset <= 1'd1;
		main_genericstandalone_rx_mmcm_reset <= 1'd1;
		main_genericstandalone_tx_init_qpll_reset0 <= 1'd0;
		main_genericstandalone_tx_init_tx_reset0 <= 1'd0;
		main_genericstandalone_tx_init_timer <= 6'd0;
		main_genericstandalone_tx_init_tick <= 1'd0;
		main_genericstandalone_rx_init_rx_reset0 <= 1'd0;
		main_genericstandalone_rx_init_drpvalue <= 16'd0;
		main_genericstandalone_rx_init_rx_pma_reset_done_r <= 1'd0;
		main_genericstandalone_cdr_lock_counter <= 13'd0;
		main_genericstandalone_cdr_locked <= 1'd0;
		main_genericstandalone_preamble_errors_status <= 32'd0;
		main_genericstandalone_crc_errors_status <= 32'd0;
		main_genericstandalone_tx_cdc_graycounter0_q <= 7'd0;
		main_genericstandalone_tx_cdc_graycounter0_q_binary <= 7'd0;
		main_genericstandalone_rx_cdc_graycounter1_q <= 7'd0;
		main_genericstandalone_rx_cdc_graycounter1_q_binary <= 7'd0;
		main_genericstandalone_sram17_status <= 32'd0;
		main_genericstandalone_sram29_storage_full <= 1'd0;
		main_genericstandalone_sram31_re <= 1'd0;
		main_genericstandalone_sram33_counter <= 11'd0;
		main_genericstandalone_slot <= 2'd0;
		main_genericstandalone_sram55_level <= 3'd0;
		main_genericstandalone_sram57_produce <= 2'd0;
		main_genericstandalone_sram58_consume <= 2'd0;
		main_genericstandalone_sram99_storage_full <= 2'd0;
		main_genericstandalone_sram101_re <= 1'd0;
		main_genericstandalone_sram102_storage_full <= 11'd0;
		main_genericstandalone_sram104_re <= 1'd0;
		main_genericstandalone_sram107_pending <= 1'd0;
		main_genericstandalone_sram116_storage_full <= 1'd0;
		main_genericstandalone_sram118_re <= 1'd0;
		main_genericstandalone_sram135_level <= 3'd0;
		main_genericstandalone_sram137_produce <= 2'd0;
		main_genericstandalone_sram138_consume <= 2'd0;
		main_genericstandalone_sram152_counter <= 11'd0;
		main_genericstandalone_last_d <= 1'd0;
		main_genericstandalone_sram0_bus_ack <= 1'd0;
		main_genericstandalone_sram1_bus_ack <= 1'd0;
		main_genericstandalone_sram2_bus_ack <= 1'd0;
		main_genericstandalone_sram3_bus_ack <= 1'd0;
		main_genericstandalone_sram4_bus_ack <= 1'd0;
		main_genericstandalone_sram5_bus_ack <= 1'd0;
		main_genericstandalone_sram6_bus_ack <= 1'd0;
		main_genericstandalone_sram7_bus_ack <= 1'd0;
		main_genericstandalone_slave_sel_r <= 8'd0;
		main_genericstandalone_kernel_cpu_storage_full <= 1'd1;
		main_genericstandalone_kernel_cpu_re <= 1'd0;
		main_genericstandalone_mailbox_i1_dat_r <= 32'd0;
		main_genericstandalone_mailbox_i1_ack <= 1'd0;
		main_genericstandalone_mailbox_i2_dat_r <= 32'd0;
		main_genericstandalone_mailbox_i2_ack <= 1'd0;
		main_genericstandalone_mailbox0 <= 32'd0;
		main_genericstandalone_mailbox1 <= 32'd0;
		main_genericstandalone_mailbox2 <= 32'd0;
		main_genericstandalone_add_identifier_storage_full <= 8'd0;
		main_genericstandalone_add_identifier_re <= 1'd0;
		main_genericstandalone_error_led_storage_full <= 1'd0;
		main_genericstandalone_error_led_re <= 1'd0;
		main_genericstandalone_rtiosyscrg_storage_full <= 1'd0;
		main_genericstandalone_rtiosyscrg_re <= 1'd0;
		main_genericstandalone_i2c_out_storage_full <= 2'd0;
		main_genericstandalone_i2c_out_re <= 1'd0;
		main_genericstandalone_i2c_oe_storage_full <= 2'd0;
		main_genericstandalone_i2c_oe_re <= 1'd0;
		main_genericstandalone_coarse_ts <= 61'd0;
		main_genericstandalone_rtio_core_storage_full <= 1'd0;
		main_genericstandalone_rtio_core_re <= 1'd0;
		main_genericstandalone_rtio_core_collision_channel_status <= 16'd0;
		main_genericstandalone_rtio_core_busy_channel_status <= 16'd0;
		main_genericstandalone_rtio_core_sequence_error_channel_status <= 16'd0;
		main_genericstandalone_rtio_core_cmd_reset <= 1'd1;
		main_genericstandalone_rtio_core_cmd_reset_phy <= 1'd1;
		main_genericstandalone_rtio_core_sed_lane_dist_minimum_coarse_timestamp <= 61'd0;
		main_genericstandalone_rtio_core_o_collision <= 1'd0;
		main_genericstandalone_rtio_core_o_busy <= 1'd0;
		main_genericstandalone_rtio_core_o_sequence_error <= 1'd0;
		main_genericstandalone_rtio_target_storage_full <= 32'd0;
		main_genericstandalone_rtio_target_re <= 1'd0;
		main_genericstandalone_rtio_o_data_storage_full <= 512'd0;
		main_genericstandalone_rtio_o_data_re <= 1'd0;
		main_genericstandalone_rtio_i_timeout_storage_full <= 64'd0;
		main_genericstandalone_rtio_i_timeout_re <= 1'd0;
		main_genericstandalone_rtio_counter_status <= 64'd0;
		main_genericstandalone_rtio_now_hi_backing <= 32'd0;
		main_genericstandalone_dma_dma_storage_full <= 33'd0;
		main_genericstandalone_dma_dma_re <= 1'd0;
		main_genericstandalone_dma_time_offset_storage_full <= 64'd0;
		main_genericstandalone_dma_time_offset_re <= 1'd0;
		main_genericstandalone_interface0_csr_bus_dat_r <= 32'd0;
		main_genericstandalone_interface0_csr_bus_ack <= 1'd0;
		main_genericstandalone_interface1_csr_bus_dat_r <= 32'd0;
		main_genericstandalone_interface1_csr_bus_ack <= 1'd0;
		main_genericstandalone_cri_con_storage_full <= 2'd0;
		main_genericstandalone_cri_con_re <= 1'd0;
		main_genericstandalone_cri_con_selected <= 1'd0;
		main_genericstandalone_interface2_csr_bus_dat_r <= 32'd0;
		main_genericstandalone_interface2_csr_bus_ack <= 1'd0;
		main_genericstandalone_mon_chan_sel_storage_full <= 6'd0;
		main_genericstandalone_mon_chan_sel_re <= 1'd0;
		main_genericstandalone_mon_probe_sel_storage_full <= 5'd0;
		main_genericstandalone_mon_probe_sel_re <= 1'd0;
		main_genericstandalone_mon_status <= 32'd0;
		main_genericstandalone_mon_bussynchronizer20_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer21_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer22_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer23_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer29_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer30_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer31_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer32_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer39_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer40_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer41_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer42_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer43_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer44_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer45_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer46_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer47_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer48_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer49_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer50_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer51_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer52_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer53_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer54_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer55_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer56_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer57_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer58_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer59_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer60_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer61_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer62_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer63_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer64_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer65_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer66_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer67_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer68_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer69_ping_o1 <= 1'd0;
		main_genericstandalone_mon_bussynchronizer70_ping_o1 <= 1'd0;
		main_genericstandalone_inj_chan_sel_storage_full <= 6'd0;
		main_genericstandalone_inj_chan_sel_re <= 1'd0;
		main_genericstandalone_inj_override_sel_storage_full <= 2'd0;
		main_genericstandalone_inj_override_sel_re <= 1'd0;
		main_genericstandalone_inj_o_sys0 <= 1'd0;
		main_genericstandalone_inj_o_sys1 <= 1'd0;
		main_genericstandalone_inj_o_sys2 <= 1'd0;
		main_genericstandalone_inj_o_sys3 <= 1'd0;
		main_genericstandalone_inj_o_sys4 <= 1'd0;
		main_genericstandalone_inj_o_sys5 <= 1'd0;
		main_genericstandalone_inj_o_sys6 <= 1'd0;
		main_genericstandalone_inj_o_sys7 <= 1'd0;
		main_genericstandalone_inj_o_sys8 <= 1'd0;
		main_genericstandalone_inj_o_sys9 <= 1'd0;
		main_genericstandalone_inj_o_sys10 <= 1'd0;
		main_genericstandalone_inj_o_sys11 <= 1'd0;
		main_genericstandalone_inj_o_sys12 <= 1'd0;
		main_genericstandalone_inj_o_sys13 <= 1'd0;
		main_genericstandalone_inj_o_sys14 <= 1'd0;
		main_genericstandalone_inj_o_sys15 <= 1'd0;
		main_genericstandalone_inj_o_sys16 <= 1'd0;
		main_genericstandalone_inj_o_sys17 <= 1'd0;
		main_genericstandalone_inj_o_sys18 <= 1'd0;
		main_genericstandalone_inj_o_sys19 <= 1'd0;
		main_genericstandalone_inj_o_sys20 <= 1'd0;
		main_genericstandalone_inj_o_sys21 <= 1'd0;
		main_genericstandalone_inj_o_sys22 <= 1'd0;
		main_genericstandalone_inj_o_sys23 <= 1'd0;
		main_genericstandalone_inj_o_sys24 <= 1'd0;
		main_genericstandalone_inj_o_sys25 <= 1'd0;
		main_genericstandalone_inj_o_sys26 <= 1'd0;
		main_genericstandalone_inj_o_sys27 <= 1'd0;
		main_genericstandalone_inj_o_sys28 <= 1'd0;
		main_genericstandalone_inj_o_sys29 <= 1'd0;
		main_genericstandalone_inj_o_sys30 <= 1'd0;
		main_genericstandalone_inj_o_sys31 <= 1'd0;
		main_genericstandalone_inj_o_sys32 <= 1'd0;
		main_genericstandalone_inj_o_sys33 <= 1'd0;
		main_genericstandalone_inj_o_sys34 <= 1'd0;
		main_genericstandalone_inj_o_sys35 <= 1'd0;
		main_genericstandalone_inj_o_sys36 <= 1'd0;
		main_genericstandalone_inj_o_sys37 <= 1'd0;
		main_genericstandalone_inj_o_sys38 <= 1'd0;
		main_genericstandalone_inj_o_sys39 <= 1'd0;
		main_genericstandalone_inj_o_sys40 <= 1'd0;
		main_genericstandalone_inj_o_sys41 <= 1'd0;
		main_genericstandalone_inj_o_sys42 <= 1'd0;
		main_genericstandalone_inj_o_sys43 <= 1'd0;
		main_genericstandalone_inj_o_sys44 <= 1'd0;
		main_genericstandalone_inj_o_sys45 <= 1'd0;
		main_genericstandalone_inj_o_sys46 <= 1'd0;
		main_genericstandalone_inj_o_sys47 <= 1'd0;
		main_genericstandalone_inj_o_sys48 <= 1'd0;
		main_genericstandalone_inj_o_sys49 <= 1'd0;
		main_genericstandalone_inj_o_sys50 <= 1'd0;
		main_genericstandalone_inj_o_sys51 <= 1'd0;
		main_genericstandalone_inj_o_sys52 <= 1'd0;
		main_genericstandalone_inj_o_sys53 <= 1'd0;
		main_genericstandalone_inj_o_sys54 <= 1'd0;
		main_genericstandalone_inj_o_sys55 <= 1'd0;
		main_genericstandalone_inj_o_sys56 <= 1'd0;
		main_genericstandalone_inj_o_sys57 <= 1'd0;
		main_genericstandalone_inj_o_sys58 <= 1'd0;
		main_genericstandalone_inj_o_sys59 <= 1'd0;
		main_genericstandalone_inj_o_sys60 <= 1'd0;
		main_genericstandalone_inj_o_sys61 <= 1'd0;
		main_genericstandalone_inj_o_sys62 <= 1'd0;
		main_genericstandalone_inj_o_sys63 <= 1'd0;
		main_genericstandalone_inj_o_sys64 <= 1'd0;
		main_genericstandalone_inj_o_sys65 <= 1'd0;
		main_genericstandalone_inj_o_sys66 <= 1'd0;
		main_genericstandalone_inj_o_sys67 <= 1'd0;
		main_genericstandalone_interface1_bus_adr <= 29'd0;
		main_genericstandalone_rtio_analyzer_enable_storage_full <= 1'd0;
		main_genericstandalone_rtio_analyzer_enable_re <= 1'd0;
		main_genericstandalone_rtio_analyzer_busy_status <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_source_stb <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_source_eop <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_source_payload_data <= 256'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_status <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_read_wait_event_r <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_just_written <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_enable_r <= 1'd0;
		main_genericstandalone_rtio_analyzer_message_encoder_stopping <= 1'd0;
		main_genericstandalone_rtio_analyzer_fifo_readable <= 1'd0;
		main_genericstandalone_rtio_analyzer_fifo_level0 <= 8'd0;
		main_genericstandalone_rtio_analyzer_fifo_produce <= 7'd0;
		main_genericstandalone_rtio_analyzer_fifo_consume <= 7'd0;
		main_genericstandalone_rtio_analyzer_fifo_transfer_count <= 6'd63;
		main_genericstandalone_rtio_analyzer_fifo_activated <= 1'd0;
		main_genericstandalone_rtio_analyzer_fifo_eop_count <= 8'd0;
		main_genericstandalone_rtio_analyzer_converter_mux <= 1'd0;
		main_genericstandalone_rtio_analyzer_dma_base_address_storage_full <= 33'd0;
		main_genericstandalone_rtio_analyzer_dma_base_address_re <= 1'd0;
		main_genericstandalone_rtio_analyzer_dma_last_address_storage_full <= 33'd0;
		main_genericstandalone_rtio_analyzer_dma_last_address_re <= 1'd0;
		main_genericstandalone_rtio_analyzer_dma_message_count <= 59'd0;
		main_genericstandalone_rtio_analyzer_enable_r <= 1'd0;
		builder_minicon_state <= 6'd0;
		builder_cache_state <= 3'd0;
		builder_a7_1000basex_gtptxinit_state <= 2'd0;
		builder_a7_1000basex_gtprxinit_state <= 4'd0;
		builder_liteethmacsramwriter_state <= 2'd0;
		builder_liteethmacsramreader_state <= 2'd0;
		builder_grant <= 1'd0;
		builder_slave_sel_r <= 5'd0;
		builder_sdram_cpulevel_arbiter_grant <= 1'd0;
		builder_sdram_native_arbiter_grant <= 2'd0;
		builder_genericstandalone_grant <= 1'd0;
		builder_genericstandalone_slave_sel_r <= 6'd0;
		builder_genericstandalone_interface0_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface1_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface2_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface3_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface4_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface5_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface6_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface7_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface8_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface9_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface10_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface11_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface12_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface13_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface14_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface15_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface16_bank_bus_dat_r <= 8'd0;
	end
	builder_xilinxmultiregimpl00 <= serial_rx;
	builder_xilinxmultiregimpl01 <= builder_xilinxmultiregimpl00;
	builder_xilinxmultiregimpl20 <= main_genericstandalone_genericstandalone_crg_o_clk_sw;
	builder_xilinxmultiregimpl21 <= builder_xilinxmultiregimpl20;
	builder_xilinxmultiregimpl100 <= main_genericstandalone_tx_init_qpll_lock0;
	builder_xilinxmultiregimpl101 <= builder_xilinxmultiregimpl100;
	builder_xilinxmultiregimpl110 <= main_genericstandalone_rx_init_rx_pma_reset_done0;
	builder_xilinxmultiregimpl111 <= builder_xilinxmultiregimpl110;
	builder_xilinxmultiregimpl120 <= main_genericstandalone_toggle_i;
	builder_xilinxmultiregimpl121 <= builder_xilinxmultiregimpl120;
	builder_xilinxmultiregimpl130 <= main_genericstandalone_ps_preamble_error_toggle_i;
	builder_xilinxmultiregimpl131 <= builder_xilinxmultiregimpl130;
	builder_xilinxmultiregimpl140 <= main_genericstandalone_ps_crc_error_toggle_i;
	builder_xilinxmultiregimpl141 <= builder_xilinxmultiregimpl140;
	builder_xilinxmultiregimpl160 <= main_genericstandalone_tx_cdc_graycounter1_q;
	builder_xilinxmultiregimpl161 <= builder_xilinxmultiregimpl160;
	builder_xilinxmultiregimpl170 <= main_genericstandalone_rx_cdc_graycounter0_q;
	builder_xilinxmultiregimpl171 <= builder_xilinxmultiregimpl170;
	builder_xilinxmultiregimpl190 <= main_genericstandalone_i2c_tstriple0_i;
	builder_xilinxmultiregimpl191 <= builder_xilinxmultiregimpl190;
	builder_xilinxmultiregimpl200 <= main_genericstandalone_i2c_tstriple1_i;
	builder_xilinxmultiregimpl201 <= builder_xilinxmultiregimpl200;
	builder_xilinxmultiregimpl220 <= main_genericstandalone_rtio_core_o_collision_sync_ps_toggle_i;
	builder_xilinxmultiregimpl221 <= builder_xilinxmultiregimpl220;
	builder_xilinxmultiregimpl240 <= main_genericstandalone_rtio_core_o_collision_sync_bxfer_data;
	builder_xilinxmultiregimpl241 <= builder_xilinxmultiregimpl240;
	builder_xilinxmultiregimpl250 <= main_genericstandalone_rtio_core_o_busy_sync_ps_toggle_i;
	builder_xilinxmultiregimpl251 <= builder_xilinxmultiregimpl250;
	builder_xilinxmultiregimpl270 <= main_genericstandalone_rtio_core_o_busy_sync_bxfer_data;
	builder_xilinxmultiregimpl271 <= builder_xilinxmultiregimpl270;
	builder_xilinxmultiregimpl280 <= main_genericstandalone_mon_bussynchronizer0_i;
	builder_xilinxmultiregimpl281 <= builder_xilinxmultiregimpl280;
	builder_xilinxmultiregimpl290 <= main_genericstandalone_mon_bussynchronizer1_i;
	builder_xilinxmultiregimpl291 <= builder_xilinxmultiregimpl290;
	builder_xilinxmultiregimpl300 <= main_genericstandalone_mon_bussynchronizer2_i;
	builder_xilinxmultiregimpl301 <= builder_xilinxmultiregimpl300;
	builder_xilinxmultiregimpl310 <= main_genericstandalone_mon_bussynchronizer3_i;
	builder_xilinxmultiregimpl311 <= builder_xilinxmultiregimpl310;
	builder_xilinxmultiregimpl320 <= main_genericstandalone_mon_bussynchronizer4_i;
	builder_xilinxmultiregimpl321 <= builder_xilinxmultiregimpl320;
	builder_xilinxmultiregimpl330 <= main_genericstandalone_mon_bussynchronizer5_i;
	builder_xilinxmultiregimpl331 <= builder_xilinxmultiregimpl330;
	builder_xilinxmultiregimpl340 <= main_genericstandalone_mon_bussynchronizer6_i;
	builder_xilinxmultiregimpl341 <= builder_xilinxmultiregimpl340;
	builder_xilinxmultiregimpl350 <= main_genericstandalone_mon_bussynchronizer7_i;
	builder_xilinxmultiregimpl351 <= builder_xilinxmultiregimpl350;
	builder_xilinxmultiregimpl360 <= main_genericstandalone_mon_bussynchronizer8_i;
	builder_xilinxmultiregimpl361 <= builder_xilinxmultiregimpl360;
	builder_xilinxmultiregimpl370 <= main_genericstandalone_mon_bussynchronizer9_i;
	builder_xilinxmultiregimpl371 <= builder_xilinxmultiregimpl370;
	builder_xilinxmultiregimpl380 <= main_genericstandalone_mon_bussynchronizer10_i;
	builder_xilinxmultiregimpl381 <= builder_xilinxmultiregimpl380;
	builder_xilinxmultiregimpl390 <= main_genericstandalone_mon_bussynchronizer11_i;
	builder_xilinxmultiregimpl391 <= builder_xilinxmultiregimpl390;
	builder_xilinxmultiregimpl400 <= main_genericstandalone_mon_bussynchronizer12_i;
	builder_xilinxmultiregimpl401 <= builder_xilinxmultiregimpl400;
	builder_xilinxmultiregimpl410 <= main_genericstandalone_mon_bussynchronizer13_i;
	builder_xilinxmultiregimpl411 <= builder_xilinxmultiregimpl410;
	builder_xilinxmultiregimpl420 <= main_genericstandalone_mon_bussynchronizer14_i;
	builder_xilinxmultiregimpl421 <= builder_xilinxmultiregimpl420;
	builder_xilinxmultiregimpl430 <= main_genericstandalone_mon_bussynchronizer15_i;
	builder_xilinxmultiregimpl431 <= builder_xilinxmultiregimpl430;
	builder_xilinxmultiregimpl440 <= main_genericstandalone_mon_bussynchronizer16_i;
	builder_xilinxmultiregimpl441 <= builder_xilinxmultiregimpl440;
	builder_xilinxmultiregimpl450 <= main_genericstandalone_mon_bussynchronizer17_i;
	builder_xilinxmultiregimpl451 <= builder_xilinxmultiregimpl450;
	builder_xilinxmultiregimpl460 <= main_genericstandalone_mon_bussynchronizer18_i;
	builder_xilinxmultiregimpl461 <= builder_xilinxmultiregimpl460;
	builder_xilinxmultiregimpl470 <= main_genericstandalone_mon_bussynchronizer19_i;
	builder_xilinxmultiregimpl471 <= builder_xilinxmultiregimpl470;
	builder_xilinxmultiregimpl480 <= main_genericstandalone_mon_bussynchronizer20_ping_toggle_i;
	builder_xilinxmultiregimpl481 <= builder_xilinxmultiregimpl480;
	builder_xilinxmultiregimpl500 <= main_genericstandalone_mon_bussynchronizer20_ibuffer;
	builder_xilinxmultiregimpl501 <= builder_xilinxmultiregimpl500;
	builder_xilinxmultiregimpl510 <= main_genericstandalone_mon_bussynchronizer21_ping_toggle_i;
	builder_xilinxmultiregimpl511 <= builder_xilinxmultiregimpl510;
	builder_xilinxmultiregimpl530 <= main_genericstandalone_mon_bussynchronizer21_ibuffer;
	builder_xilinxmultiregimpl531 <= builder_xilinxmultiregimpl530;
	builder_xilinxmultiregimpl540 <= main_genericstandalone_mon_bussynchronizer22_ping_toggle_i;
	builder_xilinxmultiregimpl541 <= builder_xilinxmultiregimpl540;
	builder_xilinxmultiregimpl560 <= main_genericstandalone_mon_bussynchronizer22_ibuffer;
	builder_xilinxmultiregimpl561 <= builder_xilinxmultiregimpl560;
	builder_xilinxmultiregimpl570 <= main_genericstandalone_mon_bussynchronizer23_ping_toggle_i;
	builder_xilinxmultiregimpl571 <= builder_xilinxmultiregimpl570;
	builder_xilinxmultiregimpl590 <= main_genericstandalone_mon_bussynchronizer23_ibuffer;
	builder_xilinxmultiregimpl591 <= builder_xilinxmultiregimpl590;
	builder_xilinxmultiregimpl600 <= main_genericstandalone_mon_bussynchronizer24_i;
	builder_xilinxmultiregimpl601 <= builder_xilinxmultiregimpl600;
	builder_xilinxmultiregimpl610 <= main_genericstandalone_mon_bussynchronizer25_i;
	builder_xilinxmultiregimpl611 <= builder_xilinxmultiregimpl610;
	builder_xilinxmultiregimpl620 <= main_genericstandalone_mon_bussynchronizer26_i;
	builder_xilinxmultiregimpl621 <= builder_xilinxmultiregimpl620;
	builder_xilinxmultiregimpl630 <= main_genericstandalone_mon_bussynchronizer27_i;
	builder_xilinxmultiregimpl631 <= builder_xilinxmultiregimpl630;
	builder_xilinxmultiregimpl640 <= main_genericstandalone_mon_bussynchronizer28_i;
	builder_xilinxmultiregimpl641 <= builder_xilinxmultiregimpl640;
	builder_xilinxmultiregimpl650 <= main_genericstandalone_mon_bussynchronizer29_ping_toggle_i;
	builder_xilinxmultiregimpl651 <= builder_xilinxmultiregimpl650;
	builder_xilinxmultiregimpl670 <= main_genericstandalone_mon_bussynchronizer29_ibuffer;
	builder_xilinxmultiregimpl671 <= builder_xilinxmultiregimpl670;
	builder_xilinxmultiregimpl680 <= main_genericstandalone_mon_bussynchronizer30_ping_toggle_i;
	builder_xilinxmultiregimpl681 <= builder_xilinxmultiregimpl680;
	builder_xilinxmultiregimpl700 <= main_genericstandalone_mon_bussynchronizer30_ibuffer;
	builder_xilinxmultiregimpl701 <= builder_xilinxmultiregimpl700;
	builder_xilinxmultiregimpl710 <= main_genericstandalone_mon_bussynchronizer31_ping_toggle_i;
	builder_xilinxmultiregimpl711 <= builder_xilinxmultiregimpl710;
	builder_xilinxmultiregimpl730 <= main_genericstandalone_mon_bussynchronizer31_ibuffer;
	builder_xilinxmultiregimpl731 <= builder_xilinxmultiregimpl730;
	builder_xilinxmultiregimpl740 <= main_genericstandalone_mon_bussynchronizer32_ping_toggle_i;
	builder_xilinxmultiregimpl741 <= builder_xilinxmultiregimpl740;
	builder_xilinxmultiregimpl760 <= main_genericstandalone_mon_bussynchronizer32_ibuffer;
	builder_xilinxmultiregimpl761 <= builder_xilinxmultiregimpl760;
	builder_xilinxmultiregimpl770 <= main_genericstandalone_mon_bussynchronizer33_i;
	builder_xilinxmultiregimpl771 <= builder_xilinxmultiregimpl770;
	builder_xilinxmultiregimpl780 <= main_genericstandalone_mon_bussynchronizer34_i;
	builder_xilinxmultiregimpl781 <= builder_xilinxmultiregimpl780;
	builder_xilinxmultiregimpl790 <= main_genericstandalone_mon_bussynchronizer35_i;
	builder_xilinxmultiregimpl791 <= builder_xilinxmultiregimpl790;
	builder_xilinxmultiregimpl800 <= main_genericstandalone_mon_bussynchronizer36_i;
	builder_xilinxmultiregimpl801 <= builder_xilinxmultiregimpl800;
	builder_xilinxmultiregimpl810 <= main_genericstandalone_mon_bussynchronizer37_i;
	builder_xilinxmultiregimpl811 <= builder_xilinxmultiregimpl810;
	builder_xilinxmultiregimpl820 <= main_genericstandalone_mon_bussynchronizer38_i;
	builder_xilinxmultiregimpl821 <= builder_xilinxmultiregimpl820;
	builder_xilinxmultiregimpl830 <= main_genericstandalone_mon_bussynchronizer39_ping_toggle_i;
	builder_xilinxmultiregimpl831 <= builder_xilinxmultiregimpl830;
	builder_xilinxmultiregimpl850 <= main_genericstandalone_mon_bussynchronizer39_ibuffer;
	builder_xilinxmultiregimpl851 <= builder_xilinxmultiregimpl850;
	builder_xilinxmultiregimpl860 <= main_genericstandalone_mon_bussynchronizer40_ping_toggle_i;
	builder_xilinxmultiregimpl861 <= builder_xilinxmultiregimpl860;
	builder_xilinxmultiregimpl880 <= main_genericstandalone_mon_bussynchronizer40_ibuffer;
	builder_xilinxmultiregimpl881 <= builder_xilinxmultiregimpl880;
	builder_xilinxmultiregimpl890 <= main_genericstandalone_mon_bussynchronizer41_ping_toggle_i;
	builder_xilinxmultiregimpl891 <= builder_xilinxmultiregimpl890;
	builder_xilinxmultiregimpl910 <= main_genericstandalone_mon_bussynchronizer41_ibuffer;
	builder_xilinxmultiregimpl911 <= builder_xilinxmultiregimpl910;
	builder_xilinxmultiregimpl920 <= main_genericstandalone_mon_bussynchronizer42_ping_toggle_i;
	builder_xilinxmultiregimpl921 <= builder_xilinxmultiregimpl920;
	builder_xilinxmultiregimpl940 <= main_genericstandalone_mon_bussynchronizer42_ibuffer;
	builder_xilinxmultiregimpl941 <= builder_xilinxmultiregimpl940;
	builder_xilinxmultiregimpl950 <= main_genericstandalone_mon_bussynchronizer43_ping_toggle_i;
	builder_xilinxmultiregimpl951 <= builder_xilinxmultiregimpl950;
	builder_xilinxmultiregimpl970 <= main_genericstandalone_mon_bussynchronizer43_ibuffer;
	builder_xilinxmultiregimpl971 <= builder_xilinxmultiregimpl970;
	builder_xilinxmultiregimpl980 <= main_genericstandalone_mon_bussynchronizer44_ping_toggle_i;
	builder_xilinxmultiregimpl981 <= builder_xilinxmultiregimpl980;
	builder_xilinxmultiregimpl1000 <= main_genericstandalone_mon_bussynchronizer44_ibuffer;
	builder_xilinxmultiregimpl1001 <= builder_xilinxmultiregimpl1000;
	builder_xilinxmultiregimpl1010 <= main_genericstandalone_mon_bussynchronizer45_ping_toggle_i;
	builder_xilinxmultiregimpl1011 <= builder_xilinxmultiregimpl1010;
	builder_xilinxmultiregimpl1030 <= main_genericstandalone_mon_bussynchronizer45_ibuffer;
	builder_xilinxmultiregimpl1031 <= builder_xilinxmultiregimpl1030;
	builder_xilinxmultiregimpl1040 <= main_genericstandalone_mon_bussynchronizer46_ping_toggle_i;
	builder_xilinxmultiregimpl1041 <= builder_xilinxmultiregimpl1040;
	builder_xilinxmultiregimpl1060 <= main_genericstandalone_mon_bussynchronizer46_ibuffer;
	builder_xilinxmultiregimpl1061 <= builder_xilinxmultiregimpl1060;
	builder_xilinxmultiregimpl1070 <= main_genericstandalone_mon_bussynchronizer47_ping_toggle_i;
	builder_xilinxmultiregimpl1071 <= builder_xilinxmultiregimpl1070;
	builder_xilinxmultiregimpl1090 <= main_genericstandalone_mon_bussynchronizer47_ibuffer;
	builder_xilinxmultiregimpl1091 <= builder_xilinxmultiregimpl1090;
	builder_xilinxmultiregimpl1100 <= main_genericstandalone_mon_bussynchronizer48_ping_toggle_i;
	builder_xilinxmultiregimpl1101 <= builder_xilinxmultiregimpl1100;
	builder_xilinxmultiregimpl1120 <= main_genericstandalone_mon_bussynchronizer48_ibuffer;
	builder_xilinxmultiregimpl1121 <= builder_xilinxmultiregimpl1120;
	builder_xilinxmultiregimpl1130 <= main_genericstandalone_mon_bussynchronizer49_ping_toggle_i;
	builder_xilinxmultiregimpl1131 <= builder_xilinxmultiregimpl1130;
	builder_xilinxmultiregimpl1150 <= main_genericstandalone_mon_bussynchronizer49_ibuffer;
	builder_xilinxmultiregimpl1151 <= builder_xilinxmultiregimpl1150;
	builder_xilinxmultiregimpl1160 <= main_genericstandalone_mon_bussynchronizer50_ping_toggle_i;
	builder_xilinxmultiregimpl1161 <= builder_xilinxmultiregimpl1160;
	builder_xilinxmultiregimpl1180 <= main_genericstandalone_mon_bussynchronizer50_ibuffer;
	builder_xilinxmultiregimpl1181 <= builder_xilinxmultiregimpl1180;
	builder_xilinxmultiregimpl1190 <= main_genericstandalone_mon_bussynchronizer51_ping_toggle_i;
	builder_xilinxmultiregimpl1191 <= builder_xilinxmultiregimpl1190;
	builder_xilinxmultiregimpl1210 <= main_genericstandalone_mon_bussynchronizer51_ibuffer;
	builder_xilinxmultiregimpl1211 <= builder_xilinxmultiregimpl1210;
	builder_xilinxmultiregimpl1220 <= main_genericstandalone_mon_bussynchronizer52_ping_toggle_i;
	builder_xilinxmultiregimpl1221 <= builder_xilinxmultiregimpl1220;
	builder_xilinxmultiregimpl1240 <= main_genericstandalone_mon_bussynchronizer52_ibuffer;
	builder_xilinxmultiregimpl1241 <= builder_xilinxmultiregimpl1240;
	builder_xilinxmultiregimpl1250 <= main_genericstandalone_mon_bussynchronizer53_ping_toggle_i;
	builder_xilinxmultiregimpl1251 <= builder_xilinxmultiregimpl1250;
	builder_xilinxmultiregimpl1270 <= main_genericstandalone_mon_bussynchronizer53_ibuffer;
	builder_xilinxmultiregimpl1271 <= builder_xilinxmultiregimpl1270;
	builder_xilinxmultiregimpl1280 <= main_genericstandalone_mon_bussynchronizer54_ping_toggle_i;
	builder_xilinxmultiregimpl1281 <= builder_xilinxmultiregimpl1280;
	builder_xilinxmultiregimpl1300 <= main_genericstandalone_mon_bussynchronizer54_ibuffer;
	builder_xilinxmultiregimpl1301 <= builder_xilinxmultiregimpl1300;
	builder_xilinxmultiregimpl1310 <= main_genericstandalone_mon_bussynchronizer55_ping_toggle_i;
	builder_xilinxmultiregimpl1311 <= builder_xilinxmultiregimpl1310;
	builder_xilinxmultiregimpl1330 <= main_genericstandalone_mon_bussynchronizer55_ibuffer;
	builder_xilinxmultiregimpl1331 <= builder_xilinxmultiregimpl1330;
	builder_xilinxmultiregimpl1340 <= main_genericstandalone_mon_bussynchronizer56_ping_toggle_i;
	builder_xilinxmultiregimpl1341 <= builder_xilinxmultiregimpl1340;
	builder_xilinxmultiregimpl1360 <= main_genericstandalone_mon_bussynchronizer56_ibuffer;
	builder_xilinxmultiregimpl1361 <= builder_xilinxmultiregimpl1360;
	builder_xilinxmultiregimpl1370 <= main_genericstandalone_mon_bussynchronizer57_ping_toggle_i;
	builder_xilinxmultiregimpl1371 <= builder_xilinxmultiregimpl1370;
	builder_xilinxmultiregimpl1390 <= main_genericstandalone_mon_bussynchronizer57_ibuffer;
	builder_xilinxmultiregimpl1391 <= builder_xilinxmultiregimpl1390;
	builder_xilinxmultiregimpl1400 <= main_genericstandalone_mon_bussynchronizer58_ping_toggle_i;
	builder_xilinxmultiregimpl1401 <= builder_xilinxmultiregimpl1400;
	builder_xilinxmultiregimpl1420 <= main_genericstandalone_mon_bussynchronizer58_ibuffer;
	builder_xilinxmultiregimpl1421 <= builder_xilinxmultiregimpl1420;
	builder_xilinxmultiregimpl1430 <= main_genericstandalone_mon_bussynchronizer59_ping_toggle_i;
	builder_xilinxmultiregimpl1431 <= builder_xilinxmultiregimpl1430;
	builder_xilinxmultiregimpl1450 <= main_genericstandalone_mon_bussynchronizer59_ibuffer;
	builder_xilinxmultiregimpl1451 <= builder_xilinxmultiregimpl1450;
	builder_xilinxmultiregimpl1460 <= main_genericstandalone_mon_bussynchronizer60_ping_toggle_i;
	builder_xilinxmultiregimpl1461 <= builder_xilinxmultiregimpl1460;
	builder_xilinxmultiregimpl1480 <= main_genericstandalone_mon_bussynchronizer60_ibuffer;
	builder_xilinxmultiregimpl1481 <= builder_xilinxmultiregimpl1480;
	builder_xilinxmultiregimpl1490 <= main_genericstandalone_mon_bussynchronizer61_ping_toggle_i;
	builder_xilinxmultiregimpl1491 <= builder_xilinxmultiregimpl1490;
	builder_xilinxmultiregimpl1510 <= main_genericstandalone_mon_bussynchronizer61_ibuffer;
	builder_xilinxmultiregimpl1511 <= builder_xilinxmultiregimpl1510;
	builder_xilinxmultiregimpl1520 <= main_genericstandalone_mon_bussynchronizer62_ping_toggle_i;
	builder_xilinxmultiregimpl1521 <= builder_xilinxmultiregimpl1520;
	builder_xilinxmultiregimpl1540 <= main_genericstandalone_mon_bussynchronizer62_ibuffer;
	builder_xilinxmultiregimpl1541 <= builder_xilinxmultiregimpl1540;
	builder_xilinxmultiregimpl1550 <= main_genericstandalone_mon_bussynchronizer63_ping_toggle_i;
	builder_xilinxmultiregimpl1551 <= builder_xilinxmultiregimpl1550;
	builder_xilinxmultiregimpl1570 <= main_genericstandalone_mon_bussynchronizer63_ibuffer;
	builder_xilinxmultiregimpl1571 <= builder_xilinxmultiregimpl1570;
	builder_xilinxmultiregimpl1580 <= main_genericstandalone_mon_bussynchronizer64_ping_toggle_i;
	builder_xilinxmultiregimpl1581 <= builder_xilinxmultiregimpl1580;
	builder_xilinxmultiregimpl1600 <= main_genericstandalone_mon_bussynchronizer64_ibuffer;
	builder_xilinxmultiregimpl1601 <= builder_xilinxmultiregimpl1600;
	builder_xilinxmultiregimpl1610 <= main_genericstandalone_mon_bussynchronizer65_ping_toggle_i;
	builder_xilinxmultiregimpl1611 <= builder_xilinxmultiregimpl1610;
	builder_xilinxmultiregimpl1630 <= main_genericstandalone_mon_bussynchronizer65_ibuffer;
	builder_xilinxmultiregimpl1631 <= builder_xilinxmultiregimpl1630;
	builder_xilinxmultiregimpl1640 <= main_genericstandalone_mon_bussynchronizer66_ping_toggle_i;
	builder_xilinxmultiregimpl1641 <= builder_xilinxmultiregimpl1640;
	builder_xilinxmultiregimpl1660 <= main_genericstandalone_mon_bussynchronizer66_ibuffer;
	builder_xilinxmultiregimpl1661 <= builder_xilinxmultiregimpl1660;
	builder_xilinxmultiregimpl1670 <= main_genericstandalone_mon_bussynchronizer67_ping_toggle_i;
	builder_xilinxmultiregimpl1671 <= builder_xilinxmultiregimpl1670;
	builder_xilinxmultiregimpl1690 <= main_genericstandalone_mon_bussynchronizer67_ibuffer;
	builder_xilinxmultiregimpl1691 <= builder_xilinxmultiregimpl1690;
	builder_xilinxmultiregimpl1700 <= main_genericstandalone_mon_bussynchronizer68_ping_toggle_i;
	builder_xilinxmultiregimpl1701 <= builder_xilinxmultiregimpl1700;
	builder_xilinxmultiregimpl1720 <= main_genericstandalone_mon_bussynchronizer68_ibuffer;
	builder_xilinxmultiregimpl1721 <= builder_xilinxmultiregimpl1720;
	builder_xilinxmultiregimpl1730 <= main_genericstandalone_mon_bussynchronizer69_ping_toggle_i;
	builder_xilinxmultiregimpl1731 <= builder_xilinxmultiregimpl1730;
	builder_xilinxmultiregimpl1750 <= main_genericstandalone_mon_bussynchronizer69_ibuffer;
	builder_xilinxmultiregimpl1751 <= builder_xilinxmultiregimpl1750;
	builder_xilinxmultiregimpl1760 <= main_genericstandalone_mon_bussynchronizer70_ping_toggle_i;
	builder_xilinxmultiregimpl1761 <= builder_xilinxmultiregimpl1760;
	builder_xilinxmultiregimpl1780 <= main_genericstandalone_mon_bussynchronizer70_ibuffer;
	builder_xilinxmultiregimpl1781 <= builder_xilinxmultiregimpl1780;
	builder_xilinxmultiregimpl1790 <= main_genericstandalone_mon_bussynchronizer71_i;
	builder_xilinxmultiregimpl1791 <= builder_xilinxmultiregimpl1790;
	builder_xilinxmultiregimpl1800 <= main_genericstandalone_mon_bussynchronizer72_i;
	builder_xilinxmultiregimpl1801 <= builder_xilinxmultiregimpl1800;
	builder_xilinxmultiregimpl1810 <= main_genericstandalone_mon_bussynchronizer73_i;
	builder_xilinxmultiregimpl1811 <= builder_xilinxmultiregimpl1810;
	builder_xilinxmultiregimpl1820 <= main_genericstandalone_mon_bussynchronizer74_i;
	builder_xilinxmultiregimpl1821 <= builder_xilinxmultiregimpl1820;
	builder_xilinxmultiregimpl1830 <= main_genericstandalone_mon_bussynchronizer75_i;
	builder_xilinxmultiregimpl1831 <= builder_xilinxmultiregimpl1830;
end

always @(posedge sys_kernel_clk) begin
	main_genericstandalone_dma_dma_enable_r <= main_genericstandalone_dma_flow_enable;
	if ((main_genericstandalone_dma_flow_enable & (~main_genericstandalone_dma_dma_enable_r))) begin
		main_genericstandalone_dma_dma_sink_payload_address <= main_genericstandalone_dma_dma_storage;
		main_genericstandalone_dma_dma_sink_eop <= 1'd0;
		main_genericstandalone_dma_dma_sink_stb <= 1'd1;
	end
	if ((main_genericstandalone_dma_dma_sink_stb & main_genericstandalone_dma_dma_sink_ack)) begin
		if (main_genericstandalone_dma_dma_sink_eop) begin
			main_genericstandalone_dma_dma_sink_stb <= 1'd0;
		end else begin
			main_genericstandalone_dma_dma_sink_payload_address <= (main_genericstandalone_dma_dma_sink_payload_address + 1'd1);
			if ((~main_genericstandalone_dma_flow_enable)) begin
				main_genericstandalone_dma_dma_sink_eop <= 1'd1;
			end
		end
	end
	if (main_genericstandalone_dma_dma_transfer_cyc_rst) begin
		main_genericstandalone_dma_dma_transfer_cyc <= 6'd63;
	end else begin
		if (main_genericstandalone_dma_dma_transfer_cyc_ce) begin
			main_genericstandalone_dma_dma_transfer_cyc <= (main_genericstandalone_dma_dma_transfer_cyc - 1'd1);
		end
	end
	if ((~main_genericstandalone_dma_fifo_recv_activated)) begin
		main_genericstandalone_dma_fifo_recv_activated <= (main_genericstandalone_dma_fifo_almost_empty & (~(main_genericstandalone_dma_fifo_do_write & main_genericstandalone_dma_fifo_sink_eop)));
	end else begin
		if ((main_genericstandalone_dma_fifo_recv_activated & (main_genericstandalone_dma_fifo_do_write & (main_genericstandalone_dma_fifo_sink_last | main_genericstandalone_dma_fifo_sink_eop)))) begin
			main_genericstandalone_dma_fifo_recv_activated <= 1'd0;
		end
	end
	if (main_genericstandalone_dma_fifo_syncfifo_re) begin
		main_genericstandalone_dma_fifo_readable <= 1'd1;
	end else begin
		if (main_genericstandalone_dma_fifo_re) begin
			main_genericstandalone_dma_fifo_readable <= 1'd0;
		end
	end
	if (((main_genericstandalone_dma_fifo_syncfifo_we & main_genericstandalone_dma_fifo_syncfifo_writable) & (~main_genericstandalone_dma_fifo_replace))) begin
		main_genericstandalone_dma_fifo_produce <= (main_genericstandalone_dma_fifo_produce + 1'd1);
	end
	if (main_genericstandalone_dma_fifo_do_read) begin
		main_genericstandalone_dma_fifo_consume <= (main_genericstandalone_dma_fifo_consume + 1'd1);
	end
	if (((main_genericstandalone_dma_fifo_syncfifo_we & main_genericstandalone_dma_fifo_syncfifo_writable) & (~main_genericstandalone_dma_fifo_replace))) begin
		if ((~main_genericstandalone_dma_fifo_do_read)) begin
			main_genericstandalone_dma_fifo_level0 <= (main_genericstandalone_dma_fifo_level0 + 1'd1);
		end
	end else begin
		if (main_genericstandalone_dma_fifo_do_read) begin
			main_genericstandalone_dma_fifo_level0 <= (main_genericstandalone_dma_fifo_level0 - 1'd1);
		end
	end
	main_genericstandalone_dma_rawslicer_level <= main_genericstandalone_dma_rawslicer_next_level;
	if (main_genericstandalone_dma_rawslicer_load_buf) begin
		case (main_genericstandalone_dma_rawslicer_level)
			1'd0: begin
				main_genericstandalone_dma_rawslicer_buf[127:0] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			1'd1: begin
				main_genericstandalone_dma_rawslicer_buf[135:8] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			2'd2: begin
				main_genericstandalone_dma_rawslicer_buf[143:16] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			2'd3: begin
				main_genericstandalone_dma_rawslicer_buf[151:24] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd4: begin
				main_genericstandalone_dma_rawslicer_buf[159:32] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd5: begin
				main_genericstandalone_dma_rawslicer_buf[167:40] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd6: begin
				main_genericstandalone_dma_rawslicer_buf[175:48] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd7: begin
				main_genericstandalone_dma_rawslicer_buf[183:56] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd8: begin
				main_genericstandalone_dma_rawslicer_buf[191:64] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd9: begin
				main_genericstandalone_dma_rawslicer_buf[199:72] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd10: begin
				main_genericstandalone_dma_rawslicer_buf[207:80] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd11: begin
				main_genericstandalone_dma_rawslicer_buf[215:88] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd12: begin
				main_genericstandalone_dma_rawslicer_buf[223:96] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd13: begin
				main_genericstandalone_dma_rawslicer_buf[231:104] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd14: begin
				main_genericstandalone_dma_rawslicer_buf[239:112] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd15: begin
				main_genericstandalone_dma_rawslicer_buf[247:120] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd16: begin
				main_genericstandalone_dma_rawslicer_buf[255:128] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd17: begin
				main_genericstandalone_dma_rawslicer_buf[263:136] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd18: begin
				main_genericstandalone_dma_rawslicer_buf[271:144] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd19: begin
				main_genericstandalone_dma_rawslicer_buf[279:152] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd20: begin
				main_genericstandalone_dma_rawslicer_buf[287:160] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd21: begin
				main_genericstandalone_dma_rawslicer_buf[295:168] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd22: begin
				main_genericstandalone_dma_rawslicer_buf[303:176] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd23: begin
				main_genericstandalone_dma_rawslicer_buf[311:184] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd24: begin
				main_genericstandalone_dma_rawslicer_buf[319:192] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd25: begin
				main_genericstandalone_dma_rawslicer_buf[327:200] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd26: begin
				main_genericstandalone_dma_rawslicer_buf[335:208] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd27: begin
				main_genericstandalone_dma_rawslicer_buf[343:216] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd28: begin
				main_genericstandalone_dma_rawslicer_buf[351:224] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd29: begin
				main_genericstandalone_dma_rawslicer_buf[359:232] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd30: begin
				main_genericstandalone_dma_rawslicer_buf[367:240] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd31: begin
				main_genericstandalone_dma_rawslicer_buf[375:248] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd32: begin
				main_genericstandalone_dma_rawslicer_buf[383:256] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd33: begin
				main_genericstandalone_dma_rawslicer_buf[391:264] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd34: begin
				main_genericstandalone_dma_rawslicer_buf[399:272] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd35: begin
				main_genericstandalone_dma_rawslicer_buf[407:280] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd36: begin
				main_genericstandalone_dma_rawslicer_buf[415:288] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd37: begin
				main_genericstandalone_dma_rawslicer_buf[423:296] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd38: begin
				main_genericstandalone_dma_rawslicer_buf[431:304] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd39: begin
				main_genericstandalone_dma_rawslicer_buf[439:312] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd40: begin
				main_genericstandalone_dma_rawslicer_buf[447:320] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd41: begin
				main_genericstandalone_dma_rawslicer_buf[455:328] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd42: begin
				main_genericstandalone_dma_rawslicer_buf[463:336] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd43: begin
				main_genericstandalone_dma_rawslicer_buf[471:344] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd44: begin
				main_genericstandalone_dma_rawslicer_buf[479:352] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd45: begin
				main_genericstandalone_dma_rawslicer_buf[487:360] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd46: begin
				main_genericstandalone_dma_rawslicer_buf[495:368] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd47: begin
				main_genericstandalone_dma_rawslicer_buf[503:376] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd48: begin
				main_genericstandalone_dma_rawslicer_buf[511:384] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd49: begin
				main_genericstandalone_dma_rawslicer_buf[519:392] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd50: begin
				main_genericstandalone_dma_rawslicer_buf[527:400] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd51: begin
				main_genericstandalone_dma_rawslicer_buf[535:408] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd52: begin
				main_genericstandalone_dma_rawslicer_buf[543:416] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd53: begin
				main_genericstandalone_dma_rawslicer_buf[551:424] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd54: begin
				main_genericstandalone_dma_rawslicer_buf[559:432] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd55: begin
				main_genericstandalone_dma_rawslicer_buf[567:440] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd56: begin
				main_genericstandalone_dma_rawslicer_buf[575:448] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd57: begin
				main_genericstandalone_dma_rawslicer_buf[583:456] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd58: begin
				main_genericstandalone_dma_rawslicer_buf[591:464] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd59: begin
				main_genericstandalone_dma_rawslicer_buf[599:472] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd60: begin
				main_genericstandalone_dma_rawslicer_buf[607:480] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd61: begin
				main_genericstandalone_dma_rawslicer_buf[615:488] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd62: begin
				main_genericstandalone_dma_rawslicer_buf[623:496] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd63: begin
				main_genericstandalone_dma_rawslicer_buf[631:504] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd64: begin
				main_genericstandalone_dma_rawslicer_buf[639:512] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd65: begin
				main_genericstandalone_dma_rawslicer_buf[647:520] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd66: begin
				main_genericstandalone_dma_rawslicer_buf[655:528] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd67: begin
				main_genericstandalone_dma_rawslicer_buf[663:536] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd68: begin
				main_genericstandalone_dma_rawslicer_buf[671:544] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd69: begin
				main_genericstandalone_dma_rawslicer_buf[679:552] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd70: begin
				main_genericstandalone_dma_rawslicer_buf[687:560] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd71: begin
				main_genericstandalone_dma_rawslicer_buf[695:568] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd72: begin
				main_genericstandalone_dma_rawslicer_buf[703:576] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd73: begin
				main_genericstandalone_dma_rawslicer_buf[711:584] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd74: begin
				main_genericstandalone_dma_rawslicer_buf[719:592] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd75: begin
				main_genericstandalone_dma_rawslicer_buf[727:600] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd76: begin
				main_genericstandalone_dma_rawslicer_buf[735:608] <= {main_genericstandalone_dma_rawslicer_sink_payload_data[7:0], main_genericstandalone_dma_rawslicer_sink_payload_data[15:8], main_genericstandalone_dma_rawslicer_sink_payload_data[23:16], main_genericstandalone_dma_rawslicer_sink_payload_data[31:24], main_genericstandalone_dma_rawslicer_sink_payload_data[39:32], main_genericstandalone_dma_rawslicer_sink_payload_data[47:40], main_genericstandalone_dma_rawslicer_sink_payload_data[55:48], main_genericstandalone_dma_rawslicer_sink_payload_data[63:56], main_genericstandalone_dma_rawslicer_sink_payload_data[71:64], main_genericstandalone_dma_rawslicer_sink_payload_data[79:72], main_genericstandalone_dma_rawslicer_sink_payload_data[87:80], main_genericstandalone_dma_rawslicer_sink_payload_data[95:88], main_genericstandalone_dma_rawslicer_sink_payload_data[103:96], main_genericstandalone_dma_rawslicer_sink_payload_data[111:104], main_genericstandalone_dma_rawslicer_sink_payload_data[119:112], main_genericstandalone_dma_rawslicer_sink_payload_data[127:120]};
			end
		endcase
	end
	if (main_genericstandalone_dma_rawslicer_shift_buf) begin
		case (main_genericstandalone_dma_rawslicer_source_consume)
			1'd0: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:0];
			end
			1'd1: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:8];
			end
			2'd2: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:16];
			end
			2'd3: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:24];
			end
			3'd4: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:32];
			end
			3'd5: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:40];
			end
			3'd6: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:48];
			end
			3'd7: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:56];
			end
			4'd8: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:64];
			end
			4'd9: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:72];
			end
			4'd10: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:80];
			end
			4'd11: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:88];
			end
			4'd12: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:96];
			end
			4'd13: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:104];
			end
			4'd14: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:112];
			end
			4'd15: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:120];
			end
			5'd16: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:128];
			end
			5'd17: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:136];
			end
			5'd18: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:144];
			end
			5'd19: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:152];
			end
			5'd20: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:160];
			end
			5'd21: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:168];
			end
			5'd22: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:176];
			end
			5'd23: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:184];
			end
			5'd24: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:192];
			end
			5'd25: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:200];
			end
			5'd26: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:208];
			end
			5'd27: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:216];
			end
			5'd28: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:224];
			end
			5'd29: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:232];
			end
			5'd30: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:240];
			end
			5'd31: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:248];
			end
			6'd32: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:256];
			end
			6'd33: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:264];
			end
			6'd34: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:272];
			end
			6'd35: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:280];
			end
			6'd36: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:288];
			end
			6'd37: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:296];
			end
			6'd38: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:304];
			end
			6'd39: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:312];
			end
			6'd40: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:320];
			end
			6'd41: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:328];
			end
			6'd42: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:336];
			end
			6'd43: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:344];
			end
			6'd44: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:352];
			end
			6'd45: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:360];
			end
			6'd46: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:368];
			end
			6'd47: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:376];
			end
			6'd48: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:384];
			end
			6'd49: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:392];
			end
			6'd50: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:400];
			end
			6'd51: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:408];
			end
			6'd52: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:416];
			end
			6'd53: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:424];
			end
			6'd54: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:432];
			end
			6'd55: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:440];
			end
			6'd56: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:448];
			end
			6'd57: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:456];
			end
			6'd58: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:464];
			end
			6'd59: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:472];
			end
			6'd60: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:480];
			end
			6'd61: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:488];
			end
			6'd62: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:496];
			end
			6'd63: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:504];
			end
			7'd64: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:512];
			end
			7'd65: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:520];
			end
			7'd66: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:528];
			end
			7'd67: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:536];
			end
			7'd68: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:544];
			end
			7'd69: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:552];
			end
			7'd70: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:560];
			end
			7'd71: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:568];
			end
			7'd72: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:576];
			end
			7'd73: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:584];
			end
			7'd74: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:592];
			end
			7'd75: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:600];
			end
			7'd76: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:608];
			end
			7'd77: begin
				main_genericstandalone_dma_rawslicer_buf <= main_genericstandalone_dma_rawslicer_buf[735:616];
			end
		endcase
	end
	builder_clockdomainsrenamer_resetinserter_state <= builder_clockdomainsrenamer_resetinserter_next_state;
	if (main_genericstandalone_dma_reset) begin
		main_genericstandalone_dma_rawslicer_buf <= 736'd0;
		main_genericstandalone_dma_rawslicer_level <= 7'd0;
		builder_clockdomainsrenamer_resetinserter_state <= 2'd0;
	end
	builder_clockdomainsrenamer_recordconverter_state <= builder_clockdomainsrenamer_recordconverter_next_state;
	if (main_genericstandalone_dma_time_offset_source_ack) begin
		main_genericstandalone_dma_time_offset_source_stb <= 1'd0;
	end
	if ((~main_genericstandalone_dma_time_offset_source_stb)) begin
		main_genericstandalone_dma_time_offset_source_payload_length <= main_genericstandalone_dma_time_offset_sink_payload_length;
		main_genericstandalone_dma_time_offset_source_payload_channel <= main_genericstandalone_dma_time_offset_sink_payload_channel;
		main_genericstandalone_dma_time_offset_source_payload_address <= main_genericstandalone_dma_time_offset_sink_payload_address;
		main_genericstandalone_dma_time_offset_source_payload_data <= main_genericstandalone_dma_time_offset_sink_payload_data;
		main_genericstandalone_dma_time_offset_source_payload_timestamp <= (main_genericstandalone_dma_time_offset_sink_payload_timestamp + main_genericstandalone_dma_time_offset_storage);
		main_genericstandalone_dma_time_offset_source_eop <= main_genericstandalone_dma_time_offset_sink_eop;
		main_genericstandalone_dma_time_offset_source_stb <= main_genericstandalone_dma_time_offset_sink_stb;
	end
	if (main_genericstandalone_dma_cri_master_underflow_trigger) begin
		main_genericstandalone_dma_cri_master_error_w <= 1'd1;
		main_genericstandalone_dma_cri_master_error_channel_status <= main_genericstandalone_dma_cri_master_sink_payload_channel;
		main_genericstandalone_dma_cri_master_error_timestamp_status <= main_genericstandalone_dma_cri_master_sink_payload_timestamp;
		main_genericstandalone_dma_cri_master_error_address_status <= main_genericstandalone_dma_cri_master_sink_payload_address;
	end
	if (main_genericstandalone_dma_cri_master_link_error_trigger) begin
		main_genericstandalone_dma_cri_master_error_w <= 2'd2;
		main_genericstandalone_dma_cri_master_error_channel_status <= main_genericstandalone_dma_cri_master_sink_payload_channel;
		main_genericstandalone_dma_cri_master_error_timestamp_status <= main_genericstandalone_dma_cri_master_sink_payload_timestamp;
		main_genericstandalone_dma_cri_master_error_address_status <= main_genericstandalone_dma_cri_master_sink_payload_address;
	end
	if (main_genericstandalone_dma_cri_master_error_re) begin
		main_genericstandalone_dma_cri_master_error_w <= 1'd0;
	end
	builder_clockdomainsrenamer_crimaster_state <= builder_clockdomainsrenamer_crimaster_next_state;
	builder_clockdomainsrenamer_fsm_state <= builder_clockdomainsrenamer_fsm_next_state;
	if (sys_kernel_rst) begin
		main_genericstandalone_dma_dma_sink_stb <= 1'd0;
		main_genericstandalone_dma_dma_sink_eop <= 1'd0;
		main_genericstandalone_dma_dma_sink_payload_address <= 29'd0;
		main_genericstandalone_dma_dma_transfer_cyc <= 6'd63;
		main_genericstandalone_dma_dma_enable_r <= 1'd0;
		main_genericstandalone_dma_fifo_readable <= 1'd0;
		main_genericstandalone_dma_fifo_level0 <= 8'd0;
		main_genericstandalone_dma_fifo_produce <= 7'd0;
		main_genericstandalone_dma_fifo_consume <= 7'd0;
		main_genericstandalone_dma_fifo_recv_activated <= 1'd0;
		main_genericstandalone_dma_rawslicer_buf <= 736'd0;
		main_genericstandalone_dma_rawslicer_level <= 7'd0;
		main_genericstandalone_dma_time_offset_source_stb <= 1'd0;
		main_genericstandalone_dma_time_offset_source_eop <= 1'd0;
		main_genericstandalone_dma_time_offset_source_payload_length <= 8'd0;
		main_genericstandalone_dma_time_offset_source_payload_channel <= 24'd0;
		main_genericstandalone_dma_time_offset_source_payload_timestamp <= 64'd0;
		main_genericstandalone_dma_time_offset_source_payload_address <= 8'd0;
		main_genericstandalone_dma_time_offset_source_payload_data <= 512'd0;
		main_genericstandalone_dma_cri_master_error_w <= 2'd0;
		main_genericstandalone_dma_cri_master_error_channel_status <= 24'd0;
		main_genericstandalone_dma_cri_master_error_timestamp_status <= 64'd0;
		main_genericstandalone_dma_cri_master_error_address_status <= 16'd0;
		builder_clockdomainsrenamer_resetinserter_state <= 2'd0;
		builder_clockdomainsrenamer_recordconverter_state <= 2'd0;
		builder_clockdomainsrenamer_crimaster_state <= 3'd0;
		builder_clockdomainsrenamer_fsm_state <= 3'd0;
	end
end

VexRiscv_IMA_wide VexRiscv_IMA_wide(
	.clk(sys_clk),
	.dBusWishbone_ACK(main_genericstandalone_genericstandalone_genericstandalone_dbus_ack),
	.dBusWishbone_DAT_MISO(main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_r),
	.dBusWishbone_ERR(main_genericstandalone_genericstandalone_genericstandalone_dbus_err),
	.externalInterruptArray(main_genericstandalone_genericstandalone_genericstandalone_interrupt),
	.externalResetVector(23'd4194304),
	.iBusWishbone_ACK(main_genericstandalone_genericstandalone_genericstandalone_ibus_ack),
	.iBusWishbone_DAT_MISO(main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_r),
	.iBusWishbone_ERR(main_genericstandalone_genericstandalone_genericstandalone_ibus_err),
	.reset(sys_rst),
	.timerInterrupt(1'd0),
	.dBusWishbone_ADR(main_genericstandalone_genericstandalone_genericstandalone_dbus_adr),
	.dBusWishbone_BTE(main_genericstandalone_genericstandalone_genericstandalone_dbus_bte),
	.dBusWishbone_CTI(main_genericstandalone_genericstandalone_genericstandalone_dbus_cti),
	.dBusWishbone_CYC(main_genericstandalone_genericstandalone_genericstandalone_dbus_cyc),
	.dBusWishbone_DAT_MOSI(main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_w),
	.dBusWishbone_SEL(main_genericstandalone_genericstandalone_genericstandalone_dbus_sel),
	.dBusWishbone_STB(main_genericstandalone_genericstandalone_genericstandalone_dbus_stb),
	.dBusWishbone_WE(main_genericstandalone_genericstandalone_genericstandalone_dbus_we),
	.iBusWishbone_ADR(main_genericstandalone_genericstandalone_genericstandalone_ibus_adr),
	.iBusWishbone_BTE(main_genericstandalone_genericstandalone_genericstandalone_ibus_bte),
	.iBusWishbone_CTI(main_genericstandalone_genericstandalone_genericstandalone_ibus_cti),
	.iBusWishbone_CYC(main_genericstandalone_genericstandalone_genericstandalone_ibus_cyc),
	.iBusWishbone_DAT_MOSI(main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_w),
	.iBusWishbone_SEL(main_genericstandalone_genericstandalone_genericstandalone_ibus_sel),
	.iBusWishbone_STB(main_genericstandalone_genericstandalone_genericstandalone_ibus_stb),
	.iBusWishbone_WE(main_genericstandalone_genericstandalone_genericstandalone_ibus_we)
);

reg [63:0] mem[0:1023];
reg [9:0] memadr;
always @(posedge sys_clk) begin : mem_write_block
	integer we_index;
	for (we_index = 0; we_index < 8; we_index = we_index + 1)
		if (main_genericstandalone_genericstandalone_genericstandalone_sram_we[we_index])
			mem[main_genericstandalone_genericstandalone_genericstandalone_sram_adr][we_index * 8 +: 8] <= main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w[we_index * 8 +: 8];
	memadr <= main_genericstandalone_genericstandalone_genericstandalone_sram_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_sram_dat_r = mem[memadr];

reg [8:0] storage[0:15];
reg [8:0] memdat;
always @(posedge sys_clk) begin : mem_write_block_1
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_we)
		storage[main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr] <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_w;
	memdat <= storage[main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin : mem_write_block_2
end

assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_r = memdat;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_dat_r = storage[main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_adr];

reg [8:0] storage_1[0:15];
reg [8:0] memdat_1;
always @(posedge sys_clk) begin : mem_write_block_3
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_we)
		storage_1[main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr] <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_w;
	memdat_1 <= storage_1[main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin : mem_write_block_4
end

assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_r = memdat_1;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_dat_r = storage_1[main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_adr];

IBUFDS_GTE2 #(
	.CLKCM_CFG("TRUE"),
	.CLKRCV_TRST("TRUE"),
	.CLKSWING_CFG(2'd3)
) IBUFDS_GTE2 (
	.CEB(1'd0),
	.I(clk125_gtp_p),
	.IB(clk125_gtp_n),
	.O(main_genericstandalone_genericstandalone_crg_clk125_buf),
	.ODIV2(main_genericstandalone_genericstandalone_crg_clk125_div2_raw)
);

BUFH BUFH(
	.I(main_genericstandalone_genericstandalone_crg_clk125_div2_raw),
	.O(main_genericstandalone_genericstandalone_crg_clk125_div2)
);

PLLE2_BASE #(
	.CLKFBOUT_MULT(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE(3'd5),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(8.0),
	.CLKOUT1_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1)
) PLLE2_BASE (
	.CLKFBIN(main_genericstandalone_genericstandalone_crg_pll_fb),
	.CLKIN1(main_genericstandalone_genericstandalone_crg_clk125_div2),
	.CLKFBOUT(main_genericstandalone_genericstandalone_crg_pll_fb),
	.CLKOUT0(main_genericstandalone_genericstandalone_crg_pll_clk200),
	.CLKOUT1(main_genericstandalone_genericstandalone_crg_pll_clk_bootstrap),
	.LOCKED(main_genericstandalone_genericstandalone_crg_pll_locked)
);

BUFG BUFG(
	.I(main_genericstandalone_genericstandalone_crg_pll_clk_bootstrap),
	.O(bootstrap_clk)
);

BUFG BUFG_1(
	.I(main_genericstandalone_genericstandalone_crg_pll_clk200),
	.O(clk200_clk)
);

IDELAYCTRL IDELAYCTRL(
	.REFCLK(clk200_clk),
	.RST(main_genericstandalone_genericstandalone_crg_ic_reset)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(1'd0),
	.D2(1'd1),
	.D3(1'd0),
	.D4(1'd1),
	.D5(1'd0),
	.D6(1'd1),
	.D7(1'd0),
	.D8(1'd1),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_sd_clk_se)
);

OBUFDS OBUFDS(
	.I(main_genericstandalone_genericstandalone_ddrphy_sd_clk_se),
	.O(ddram_clk_p),
	.OB(ddram_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_1 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[0]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[0]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[0]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[0]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[0]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[0]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[1]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[1]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[1]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[1]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[1]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[1]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[1]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_3 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[2]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[2]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[2]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[2]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[2]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[2]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_4 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[3]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[3]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[3]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[3]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[3]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[3]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[3]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_5 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[4]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[4]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[4]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[4]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[4]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[4]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[4]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[4])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_6 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[5]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[5]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[5]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[5]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[5]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[5]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[5]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[5])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_7 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[6]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[6]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[6]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[6]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[6]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[6]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[6]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[6])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_8 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[7]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[7]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[7]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[7]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[7]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[7]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[7]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[7])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_9 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[8]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[8]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[8]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[8]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[8]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[8]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[8]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[8])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_10 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[9]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[9]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[9]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[9]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[9]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[9]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[9]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[9])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_11 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[10]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[10]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[10]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[10]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[10]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[10]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[10]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[10])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_12 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[11]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[11]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[11]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[11]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[11]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[11]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[11]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[11])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_13 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[12]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[12]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[12]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[12]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[12]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[12]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[12]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[12])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_14 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[13]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[13]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[13]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[13]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[13]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[13]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[13]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[13])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_15 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[14]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[14]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[14]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[14]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[14]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[14]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[14]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[14]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[14])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_16 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[0]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[0]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[0]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[0]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[0]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[0]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_17 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[1]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[1]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[1]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[1]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[1]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[1]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[1]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_18 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[2]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[2]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[2]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[2]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[2]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[2]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_19 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_ras_n),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_ras_n),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_ras_n),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_ras_n),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_ras_n),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_ras_n),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_ras_n),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_ras_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ras_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_20 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cas_n),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cas_n),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cas_n),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cas_n),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cas_n),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cas_n),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cas_n),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cas_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cas_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_21 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_we_n),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_we_n),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_we_n),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_we_n),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_we_n),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_we_n),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_we_n),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_we_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_we_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_22 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cke),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cke),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cke),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cke),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cke),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cke),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cke),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cke),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cke)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_23 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_odt),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_odt),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_odt),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_odt),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_odt),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_odt),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_odt),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_odt),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_odt)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_24 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_reset_n),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_reset_n),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_reset_n),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_reset_n),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_reset_n),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_reset_n),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_reset_n),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_reset_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_reset_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_25 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask[2]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask[0]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask[2]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask[0]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask[2]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask[0]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_26 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dqs0),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dqs_t0)
);

OBUFTDS OBUFTDS(
	.I(main_genericstandalone_genericstandalone_ddrphy_dqs0),
	.T(main_genericstandalone_genericstandalone_ddrphy_dqs_t0),
	.O(ddram_dqs_p[0]),
	.OB(ddram_dqs_n[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_27 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask[1]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask[3]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask[1]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask[3]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask[1]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask[3]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask[1]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_28 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dqs1),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dqs_t1)
);

OBUFTDS OBUFTDS_1(
	.I(main_genericstandalone_genericstandalone_ddrphy_dqs1),
	.T(main_genericstandalone_genericstandalone_ddrphy_dqs_t1),
	.O(ddram_dqs_p[1]),
	.OB(ddram_dqs_n[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_29 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[16]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[0]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[16]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[0]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[16]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[0]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[16]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o0),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed0),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[16]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[0]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[16]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[0]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[16]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[0]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[16]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay0),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed0)
);

IOBUF IOBUF(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o0),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t0),
	.IO(ddram_dq[0]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_30 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[1]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[17]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[1]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[17]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[1]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[17]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[1]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[17]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o1),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t1)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_1 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed1),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[17]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[1]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[17]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[1]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[17]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[1]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[17]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[1])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_1 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay1),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed1)
);

IOBUF IOBUF_1(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o1),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t1),
	.IO(ddram_dq[1]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_31 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[2]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[18]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[18]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[2]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[18]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[2]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[18]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o2),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t2)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_2 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed2),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[18]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[2]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[18]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[2]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[18]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[2]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[18]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[2])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_2 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay2),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed2)
);

IOBUF IOBUF_2(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o2),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t2),
	.IO(ddram_dq[2]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_32 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[3]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[19]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[3]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[19]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[3]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[19]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[3]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[19]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o3),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t3)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_3 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed3),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[19]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[3]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[19]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[3]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[19]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[3]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[19]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[3])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_3 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay3),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed3)
);

IOBUF IOBUF_3(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o3),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t3),
	.IO(ddram_dq[3]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_33 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[4]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[20]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[4]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[20]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[4]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[20]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[4]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[20]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o4),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t4)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_4 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed4),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[20]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[4]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[20]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[4]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[20]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[4]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[20]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[4])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_4 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay4),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed4)
);

IOBUF IOBUF_4(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o4),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t4),
	.IO(ddram_dq[4]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_34 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[5]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[21]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[5]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[21]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[5]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[21]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[5]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[21]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o5),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t5)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_5 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed5),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[21]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[5]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[21]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[5]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[21]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[5]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[21]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[5])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_5 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay5),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed5)
);

IOBUF IOBUF_5(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o5),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t5),
	.IO(ddram_dq[5]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_35 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[6]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[22]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[6]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[22]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[6]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[22]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[6]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[22]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o6),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t6)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_6 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed6),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[22]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[6]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[22]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[6]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[22]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[6]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[22]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[6])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_6 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay6),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed6)
);

IOBUF IOBUF_6(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o6),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t6),
	.IO(ddram_dq[6]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_36 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[7]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[23]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[7]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[23]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[7]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[23]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[7]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[23]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o7),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t7)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_7 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed7),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[23]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[7]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[23]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[7]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[23]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[7]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[23]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[7])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_7 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay7),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed7)
);

IOBUF IOBUF_7(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o7),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t7),
	.IO(ddram_dq[7]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_37 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[8]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[24]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[8]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[24]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[8]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[24]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[8]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[24]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o8),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t8)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_8 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed8),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[24]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[8]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[24]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[8]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[24]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[8]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[24]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[8])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_8 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay8),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed8)
);

IOBUF IOBUF_8(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o8),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t8),
	.IO(ddram_dq[8]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay8)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_38 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[9]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[25]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[9]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[25]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[9]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[25]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[9]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[25]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o9),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t9)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_9 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed9),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[25]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[9]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[25]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[9]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[25]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[9]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[25]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[9])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_9 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay9),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed9)
);

IOBUF IOBUF_9(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o9),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t9),
	.IO(ddram_dq[9]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay9)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_39 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[10]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[26]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[10]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[26]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[10]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[26]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[10]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[26]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o10),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t10)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_10 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed10),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[26]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[10]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[26]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[10]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[26]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[10]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[26]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[10])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_10 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay10),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed10)
);

IOBUF IOBUF_10(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o10),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t10),
	.IO(ddram_dq[10]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay10)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_40 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[11]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[27]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[11]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[27]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[11]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[27]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[11]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[27]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o11),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t11)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_11 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed11),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[27]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[11]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[27]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[11]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[27]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[11]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[27]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[11])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_11 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay11),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed11)
);

IOBUF IOBUF_11(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o11),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t11),
	.IO(ddram_dq[11]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay11)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_41 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[12]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[28]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[12]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[28]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[12]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[28]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[12]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[28]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o12),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t12)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_12 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed12),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[28]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[12]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[28]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[12]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[28]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[12]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[28]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[12])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_12 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay12),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed12)
);

IOBUF IOBUF_12(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o12),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t12),
	.IO(ddram_dq[12]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay12)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_42 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[13]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[29]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[13]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[29]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[13]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[29]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[13]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[29]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o13),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t13)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_13 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed13),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[29]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[13]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[29]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[13]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[29]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[13]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[29]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[13])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_13 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay13),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed13)
);

IOBUF IOBUF_13(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o13),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t13),
	.IO(ddram_dq[13]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay13)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_43 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[14]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[30]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[14]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[30]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[14]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[30]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[14]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[30]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o14),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t14)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_14 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed14),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[30]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[14]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[30]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[14]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[30]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[14]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[30]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[14])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_14 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay14),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed14)
);

IOBUF IOBUF_14(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o14),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t14),
	.IO(ddram_dq[14]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay14)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_44 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[15]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[31]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[15]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[31]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[15]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[31]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[15]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[31]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o15),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t15)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_15 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed15),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[31]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[15]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[31]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[15]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[31]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[15]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[31]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[15])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_15 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay15),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed15)
);

IOBUF IOBUF_15(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o15),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t15),
	.IO(ddram_dq[15]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay15)
);

reg [511:0] data_mem[0:2047];
reg [10:0] memadr_1;
always @(posedge sys_clk) begin : mem_write_block_5
	integer we_index_1;
	for (we_index_1 = 0; we_index_1 < 64; we_index_1 = we_index_1 + 1)
		if (main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_we[we_index_1])
			data_mem[main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_adr][we_index_1 * 8 +: 8] <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_w[we_index_1 * 8 +: 8];
	memadr_1 <= main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_cache_data_port_dat_r = data_mem[memadr_1];

reg [16:0] tag_mem[0:2047];
reg [10:0] memadr_2;
always @(posedge sys_clk) begin : mem_write_block_6
	if (main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_we)
		tag_mem[main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_dat_w;
	memadr_2 <= main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_cache_tag_port_dat_r = tag_mem[memadr_2];

STARTUPE2 STARTUPE2(
	.CLK(1'd0),
	.GSR(1'd0),
	.GTS(1'd0),
	.KEYCLEARB(1'd0),
	.PACK(1'd0),
	.USRCCLKO(main_genericstandalone_genericstandalone_clk),
	.USRCCLKTS(1'd0),
	.USRDONEO(1'd1),
	.USRDONETS(1'd1)
);

assign spiflash2x_dq = main_genericstandalone_genericstandalone_spiflash_oe ? main_genericstandalone_genericstandalone_spiflash_o : 2'bz;
assign main_genericstandalone_genericstandalone_spiflash_i0 = spiflash2x_dq;

BUFHCE BUFHCE(
	.CE(main_genericstandalone_genericstandalone_icap_counter_rst),
	.I(sys_clk),
	.O(icap_clk)
);

ICAPE2 #(
	.ICAP_WIDTH("X32")
) ICAPE2 (
	.CLK(icap_clk),
	.CSIB(main_genericstandalone_genericstandalone_icap_icap_csib),
	.I(main_genericstandalone_genericstandalone_icap_icap_i),
	.RDWRB(main_genericstandalone_genericstandalone_icap_icap_rdwrb)
);

GTPE2_COMMON #(
	.PLL0_FBDIV(3'd4),
	.PLL0_FBDIV_45(3'd5),
	.PLL0_REFCLK_DIV(1'd1)
) GTPE2_COMMON (
	.BGBYPASSB(1'd1),
	.BGMONITORENB(1'd1),
	.BGPDB(1'd1),
	.BGRCALOVRD(5'd31),
	.GTREFCLK0(main_genericstandalone_genericstandalone_crg_clk125_buf),
	.GTREFCLK1(1'd0),
	.PLL0LOCKEN(1'd1),
	.PLL0PD(1'd0),
	.PLL0REFCLKSEL(1'd1),
	.PLL0RESET(main_genericstandalone_genericstandalone_qpll_reset),
	.PLL1PD(1'd1),
	.RCALENB(1'd1),
	.PLL0LOCK(main_genericstandalone_genericstandalone_qpll_lock),
	.PLL0OUTCLK(main_genericstandalone_genericstandalone_qpll_clk),
	.PLL0OUTREFCLK(main_genericstandalone_genericstandalone_qpll_refclk)
);

GTPE2_CHANNEL #(
	.ACJTAG_DEBUG_MODE(1'd0),
	.ACJTAG_MODE(1'd0),
	.ACJTAG_RESET(1'd0),
	.ADAPT_CFG0(1'd0),
	.ALIGN_COMMA_DOUBLE("FALSE"),
	.ALIGN_COMMA_ENABLE(10'd1023),
	.ALIGN_COMMA_WORD(1'd1),
	.ALIGN_MCOMMA_DET("TRUE"),
	.ALIGN_MCOMMA_VALUE(10'd643),
	.ALIGN_PCOMMA_DET("TRUE"),
	.ALIGN_PCOMMA_VALUE(9'd380),
	.CBCC_DATA_SOURCE_SEL("ENCODED"),
	.CFOK_CFG(43'd5016522067584),
	.CFOK_CFG2(6'd32),
	.CFOK_CFG3(6'd32),
	.CFOK_CFG4(1'd0),
	.CFOK_CFG5(1'd0),
	.CFOK_CFG6(1'd0),
	.CHAN_BOND_KEEP_ALIGN("FALSE"),
	.CHAN_BOND_MAX_SKEW(1'd1),
	.CHAN_BOND_SEQ_1_1(1'd0),
	.CHAN_BOND_SEQ_1_2(1'd0),
	.CHAN_BOND_SEQ_1_3(1'd0),
	.CHAN_BOND_SEQ_1_4(1'd0),
	.CHAN_BOND_SEQ_1_ENABLE(4'd15),
	.CHAN_BOND_SEQ_2_1(1'd0),
	.CHAN_BOND_SEQ_2_2(1'd0),
	.CHAN_BOND_SEQ_2_3(1'd0),
	.CHAN_BOND_SEQ_2_4(1'd0),
	.CHAN_BOND_SEQ_2_ENABLE(4'd15),
	.CHAN_BOND_SEQ_2_USE("FALSE"),
	.CHAN_BOND_SEQ_LEN(1'd1),
	.CLK_COMMON_SWING(1'd0),
	.CLK_CORRECT_USE("FALSE"),
	.CLK_COR_KEEP_IDLE("FALSE"),
	.CLK_COR_MAX_LAT(4'd9),
	.CLK_COR_MIN_LAT(3'd7),
	.CLK_COR_PRECEDENCE("TRUE"),
	.CLK_COR_REPEAT_WAIT(1'd0),
	.CLK_COR_SEQ_1_1(9'd256),
	.CLK_COR_SEQ_1_2(1'd0),
	.CLK_COR_SEQ_1_3(1'd0),
	.CLK_COR_SEQ_1_4(1'd0),
	.CLK_COR_SEQ_1_ENABLE(4'd15),
	.CLK_COR_SEQ_2_1(9'd256),
	.CLK_COR_SEQ_2_2(1'd0),
	.CLK_COR_SEQ_2_3(1'd0),
	.CLK_COR_SEQ_2_4(1'd0),
	.CLK_COR_SEQ_2_ENABLE(4'd15),
	.CLK_COR_SEQ_2_USE("FALSE"),
	.CLK_COR_SEQ_LEN(1'd1),
	.DEC_MCOMMA_DETECT("FALSE"),
	.DEC_PCOMMA_DETECT("FALSE"),
	.DEC_VALID_COMMA_ONLY("FALSE"),
	.DMONITOR_CFG(12'd2560),
	.ES_CLK_PHASE_SEL(1'd0),
	.ES_CONTROL(1'd0),
	.ES_ERRDET_EN("FALSE"),
	.ES_EYE_SCAN_EN("FALSE"),
	.ES_HORZ_OFFSET(5'd16),
	.ES_PMA_CFG(1'd0),
	.ES_PRESCALE(1'd0),
	.ES_QUALIFIER(1'd0),
	.ES_QUAL_MASK(1'd0),
	.ES_SDATA_MASK(1'd0),
	.ES_VERT_OFFSET(1'd0),
	.FTS_DESKEW_SEQ_ENABLE(4'd15),
	.FTS_LANE_DESKEW_CFG(4'd15),
	.FTS_LANE_DESKEW_EN("FALSE"),
	.GEARBOX_MODE(1'd0),
	.LOOPBACK_CFG(1'd0),
	.OUTREFCLK_SEL_INV(2'd3),
	.PCS_PCIE_EN("FALSE"),
	.PCS_RSVD_ATTR(1'd0),
	.PD_TRANS_TIME_FROM_P2(6'd60),
	.PD_TRANS_TIME_NONE_P2(6'd60),
	.PD_TRANS_TIME_TO_P2(7'd100),
	.PMA_LOOPBACK_CFG(1'd0),
	.PMA_RSV(10'd819),
	.PMA_RSV2(14'd8256),
	.PMA_RSV3(1'd0),
	.PMA_RSV4(1'd0),
	.PMA_RSV5(1'd0),
	.PMA_RSV6(1'd0),
	.PMA_RSV7(1'd0),
	.RXBUFRESET_TIME(1'd1),
	.RXBUF_ADDR_MODE("FAST"),
	.RXBUF_EIDLE_HI_CNT(4'd8),
	.RXBUF_EIDLE_LO_CNT(1'd0),
	.RXBUF_EN("TRUE"),
	.RXBUF_RESET_ON_CB_CHANGE("TRUE"),
	.RXBUF_RESET_ON_COMMAALIGN("FALSE"),
	.RXBUF_RESET_ON_EIDLE("FALSE"),
	.RXBUF_RESET_ON_RATE_CHANGE("TRUE"),
	.RXBUF_THRESH_OVFLW(6'd61),
	.RXBUF_THRESH_OVRD("FALSE"),
	.RXBUF_THRESH_UNDFLW(3'd4),
	.RXCDRFREQRESET_TIME(1'd1),
	.RXCDRPHRESET_TIME(1'd1),
	.RXCDR_CFG(69'd314170556264376963088),
	.RXCDR_FR_RESET_ON_EIDLE(1'd0),
	.RXCDR_HOLD_DURING_EIDLE(1'd0),
	.RXCDR_LOCK_CFG(4'd9),
	.RXCDR_PH_RESET_ON_EIDLE(1'd0),
	.RXDLY_CFG(5'd31),
	.RXDLY_LCFG(6'd48),
	.RXDLY_TAP_CFG(1'd0),
	.RXGEARBOX_EN("FALSE"),
	.RXISCANRESET_TIME(1'd1),
	.RXLPMRESET_TIME(4'd15),
	.RXLPM_BIAS_STARTUP_DISABLE(1'd0),
	.RXLPM_CFG(3'd6),
	.RXLPM_CFG1(1'd0),
	.RXLPM_CM_CFG(1'd0),
	.RXLPM_GC_CFG(9'd482),
	.RXLPM_GC_CFG2(1'd1),
	.RXLPM_HF_CFG(10'd1008),
	.RXLPM_HF_CFG2(4'd10),
	.RXLPM_HF_CFG3(1'd0),
	.RXLPM_HOLD_DURING_EIDLE(1'd0),
	.RXLPM_INCM_CFG(1'd0),
	.RXLPM_IPCM_CFG(1'd1),
	.RXLPM_LF_CFG(10'd1008),
	.RXLPM_LF_CFG2(4'd10),
	.RXLPM_OSINT_CFG(3'd4),
	.RXOOB_CFG(3'd6),
	.RXOOB_CLK_CFG("PMA"),
	.RXOSCALRESET_TIME(2'd3),
	.RXOSCALRESET_TIMEOUT(1'd0),
	.RXOUT_DIV(3'd4),
	.RXPCSRESET_TIME(1'd1),
	.RXPHDLY_CFG(20'd540704),
	.RXPH_CFG(24'd12582914),
	.RXPH_MONITOR_SEL(1'd0),
	.RXPI_CFG0(1'd0),
	.RXPI_CFG1(1'd1),
	.RXPI_CFG2(1'd1),
	.RXPMARESET_TIME(2'd3),
	.RXPRBS_ERR_LOOPBACK(1'd0),
	.RXSLIDE_AUTO_WAIT(3'd7),
	.RXSLIDE_MODE("OFF"),
	.RXSYNC_MULTILANE(1'd0),
	.RXSYNC_OVRD(1'd0),
	.RXSYNC_SKIP_DA(1'd0),
	.RX_BIAS_CFG(12'd3891),
	.RX_BUFFER_CFG(1'd0),
	.RX_CLK25_DIV(3'd5),
	.RX_CLKMUX_EN(1'd1),
	.RX_CM_SEL(1'd1),
	.RX_CM_TRIM(1'd0),
	.RX_DATA_WIDTH(5'd20),
	.RX_DDI_SEL(1'd0),
	.RX_DEBUG_CFG(1'd0),
	.RX_DEFER_RESET_BUF_EN("TRUE"),
	.RX_DISPERR_SEQ_MATCH("FALSE"),
	.RX_OS_CFG(8'd128),
	.RX_SIG_VALID_DLY(4'd10),
	.RX_XCLK_SEL("RXREC"),
	.SAS_MAX_COM(7'd64),
	.SAS_MIN_COM(6'd36),
	.SATA_BURST_SEQ_LEN(3'd5),
	.SATA_BURST_VAL(3'd4),
	.SATA_EIDLE_VAL(3'd4),
	.SATA_MAX_BURST(4'd8),
	.SATA_MAX_INIT(5'd21),
	.SATA_MAX_WAKE(3'd7),
	.SATA_MIN_BURST(3'd4),
	.SATA_MIN_INIT(4'd12),
	.SATA_MIN_WAKE(3'd4),
	.SATA_PLL_CFG("VCO_3000MHZ"),
	.SHOW_REALIGN_COMMA("TRUE"),
	.SIM_RECEIVER_DETECT_PASS("TRUE"),
	.SIM_RESET_SPEEDUP("FALSE"),
	.SIM_TX_EIDLE_DRIVE_LEVEL("X"),
	.SIM_VERSION("2.0"),
	.TERM_RCAL_CFG(15'd16912),
	.TERM_RCAL_OVRD(1'd0),
	.TRANS_TIME_RATE(4'd14),
	.TST_RSV(1'd0),
	.TXBUF_EN("TRUE"),
	.TXBUF_RESET_ON_RATE_CHANGE("TRUE"),
	.TXDLY_CFG(5'd31),
	.TXDLY_LCFG(6'd48),
	.TXDLY_TAP_CFG(1'd0),
	.TXGEARBOX_EN("FALSE"),
	.TXOOB_CFG(1'd0),
	.TXOUT_DIV(3'd4),
	.TXPCSRESET_TIME(1'd1),
	.TXPHDLY_CFG(20'd540704),
	.TXPH_CFG(11'd1920),
	.TXPH_MONITOR_SEL(1'd0),
	.TXPI_CFG0(1'd0),
	.TXPI_CFG1(1'd0),
	.TXPI_CFG2(1'd0),
	.TXPI_CFG3(1'd0),
	.TXPI_CFG4(1'd0),
	.TXPI_CFG5(1'd0),
	.TXPI_GREY_SEL(1'd0),
	.TXPI_INVSTROBE_SEL(1'd0),
	.TXPI_PPMCLK_SEL("TXUSRCLK2"),
	.TXPI_PPM_CFG(1'd0),
	.TXPI_SYNFREQ_PPM(1'd1),
	.TXPMARESET_TIME(1'd1),
	.TXSYNC_MULTILANE(1'd0),
	.TXSYNC_OVRD(1'd0),
	.TXSYNC_SKIP_DA(1'd0),
	.TX_CLK25_DIV(3'd5),
	.TX_CLKMUX_EN(1'd1),
	.TX_DATA_WIDTH(5'd20),
	.TX_DEEMPH0(1'd0),
	.TX_DEEMPH1(1'd0),
	.TX_DRIVE_MODE("DIRECT"),
	.TX_EIDLE_ASSERT_DELAY(3'd6),
	.TX_EIDLE_DEASSERT_DELAY(3'd4),
	.TX_LOOPBACK_DRIVE_HIZ("FALSE"),
	.TX_MAINCURSOR_SEL(1'd0),
	.TX_MARGIN_FULL_0(7'd78),
	.TX_MARGIN_FULL_1(7'd73),
	.TX_MARGIN_FULL_2(7'd69),
	.TX_MARGIN_FULL_3(7'd66),
	.TX_MARGIN_FULL_4(7'd64),
	.TX_MARGIN_LOW_0(7'd70),
	.TX_MARGIN_LOW_1(7'd68),
	.TX_MARGIN_LOW_2(7'd66),
	.TX_MARGIN_LOW_3(7'd64),
	.TX_MARGIN_LOW_4(7'd64),
	.TX_PREDRIVER_MODE(1'd0),
	.TX_RXDETECT_CFG(13'd6194),
	.TX_RXDETECT_REF(3'd4),
	.TX_XCLK_SEL("TXOUT"),
	.UCODEER_CLR(1'd0),
	.USE_PCS_CLK_PHASE_SEL(1'd0)
) GTPE2_CHANNEL (
	.CFGRESET(1'd0),
	.CLKRSVD0(1'd0),
	.CLKRSVD1(1'd0),
	.DMONFIFORESET(1'd0),
	.DMONITORCLK(1'd0),
	.DRPADDR(main_genericstandalone_drpaddr),
	.DRPCLK(sys_clk),
	.DRPDI(main_genericstandalone_drpdi),
	.DRPEN(main_genericstandalone_drpen),
	.DRPWE(main_genericstandalone_drpwe),
	.EYESCANMODE(1'd0),
	.EYESCANRESET(1'd0),
	.EYESCANTRIGGER(1'd0),
	.GTPRXN(sfp_rxn),
	.GTPRXP(sfp_rxp),
	.GTRESETSEL(1'd0),
	.GTRSVD(1'd0),
	.GTRXRESET(main_genericstandalone_rx_reset),
	.GTTXRESET(main_genericstandalone_tx_reset),
	.LOOPBACK(1'd0),
	.PCSRSVDIN(1'd0),
	.PLL0CLK(main_genericstandalone_genericstandalone_qpll_clk),
	.PLL0REFCLK(main_genericstandalone_genericstandalone_qpll_refclk),
	.PLL1CLK(1'd0),
	.PLL1REFCLK(1'd0),
	.PMARSVDIN0(1'd0),
	.PMARSVDIN1(1'd0),
	.PMARSVDIN2(1'd0),
	.PMARSVDIN3(1'd0),
	.PMARSVDIN4(1'd0),
	.RESETOVRD(1'd0),
	.RX8B10BEN(1'd0),
	.RXADAPTSELTEST(1'd0),
	.RXBUFRESET(1'd0),
	.RXCDRFREQRESET(1'd0),
	.RXCDRHOLD(1'd0),
	.RXCDROVRDEN(1'd0),
	.RXCDRRESET(1'd0),
	.RXCDRRESETRSV(1'd0),
	.RXCHBONDEN(1'd0),
	.RXCHBONDI(1'd0),
	.RXCHBONDLEVEL(1'd0),
	.RXCHBONDMASTER(1'd0),
	.RXCHBONDSLAVE(1'd0),
	.RXCOMMADETEN(1'd0),
	.RXDDIEN(1'd0),
	.RXDFEXYDEN(1'd0),
	.RXDLYBYPASS(1'd1),
	.RXDLYEN(1'd0),
	.RXDLYOVRDEN(1'd0),
	.RXDLYSRESET(1'd0),
	.RXELECIDLEMODE(2'd3),
	.RXGEARBOXSLIP(1'd0),
	.RXLPMHFHOLD(1'd0),
	.RXLPMHFOVRDEN(1'd0),
	.RXLPMLFHOLD(1'd0),
	.RXLPMLFOVRDEN(1'd0),
	.RXLPMOSINTNTRLEN(1'd0),
	.RXLPMRESET(1'd0),
	.RXMCOMMAALIGNEN(1'd0),
	.RXOOBRESET(1'd0),
	.RXOSCALRESET(1'd0),
	.RXOSHOLD(1'd0),
	.RXOSINTCFG(2'd2),
	.RXOSINTEN(1'd1),
	.RXOSINTHOLD(1'd0),
	.RXOSINTID0(1'd0),
	.RXOSINTNTRLEN(1'd0),
	.RXOSINTOVRDEN(1'd0),
	.RXOSINTPD(1'd0),
	.RXOSINTSTROBE(1'd0),
	.RXOSINTTESTOVRDEN(1'd0),
	.RXOSOVRDEN(1'd0),
	.RXOUTCLKSEL(2'd2),
	.RXPCOMMAALIGNEN(1'd0),
	.RXPCSRESET(1'd0),
	.RXPD(1'd0),
	.RXPHALIGN(1'd0),
	.RXPHALIGNEN(1'd0),
	.RXPHDLYPD(1'd0),
	.RXPHDLYRESET(1'd0),
	.RXPHOVRDEN(1'd0),
	.RXPMARESET(1'd0),
	.RXPOLARITY(1'd0),
	.RXPRBSCNTRESET(1'd0),
	.RXPRBSSEL(1'd0),
	.RXRATE(1'd0),
	.RXRATEMODE(1'd0),
	.RXSLIDE(1'd0),
	.RXSYNCALLIN(1'd0),
	.RXSYNCIN(1'd0),
	.RXSYNCMODE(1'd0),
	.RXSYSCLKSEL(1'd0),
	.RXUSERRDY(main_genericstandalone_rx_mmcm_locked),
	.RXUSRCLK(eth_rx_half_clk),
	.RXUSRCLK2(eth_rx_half_clk),
	.SETERRSTATUS(1'd0),
	.SIGVALIDCLK(1'd0),
	.TSTIN(20'd1048575),
	.TX8B10BBYPASS(1'd0),
	.TX8B10BEN(1'd0),
	.TXBUFDIFFCTRL(3'd4),
	.TXCHARDISPMODE({main_genericstandalone_tx_data0[19], main_genericstandalone_tx_data0[9]}),
	.TXCHARDISPVAL({main_genericstandalone_tx_data0[18], main_genericstandalone_tx_data0[8]}),
	.TXCHARISK(1'd0),
	.TXCOMINIT(1'd0),
	.TXCOMSAS(1'd0),
	.TXCOMWAKE(1'd0),
	.TXDATA({main_genericstandalone_tx_data0[17:10], main_genericstandalone_tx_data0[7:0]}),
	.TXDEEMPH(1'd0),
	.TXDETECTRX(1'd0),
	.TXDIFFCTRL(4'd8),
	.TXDIFFPD(1'd0),
	.TXDLYBYPASS(1'd1),
	.TXDLYEN(1'd0),
	.TXDLYHOLD(1'd0),
	.TXDLYOVRDEN(1'd0),
	.TXDLYSRESET(1'd0),
	.TXDLYUPDOWN(1'd0),
	.TXELECIDLE(1'd0),
	.TXHEADER(1'd0),
	.TXINHIBIT(1'd0),
	.TXMAINCURSOR(1'd0),
	.TXMARGIN(1'd0),
	.TXOUTCLKSEL(2'd2),
	.TXPCSRESET(1'd0),
	.TXPD(1'd0),
	.TXPDELECIDLEMODE(1'd0),
	.TXPHALIGN(1'd0),
	.TXPHALIGNEN(1'd0),
	.TXPHDLYPD(1'd0),
	.TXPHDLYRESET(1'd0),
	.TXPHDLYTSTCLK(1'd0),
	.TXPHINIT(1'd0),
	.TXPHOVRDEN(1'd0),
	.TXPIPPMEN(1'd0),
	.TXPIPPMOVRDEN(1'd0),
	.TXPIPPMPD(1'd0),
	.TXPIPPMSEL(1'd1),
	.TXPIPPMSTEPSIZE(1'd0),
	.TXPISOPD(1'd0),
	.TXPMARESET(1'd0),
	.TXPOLARITY(1'd0),
	.TXPOSTCURSOR(1'd0),
	.TXPOSTCURSORINV(1'd0),
	.TXPRBSFORCEERR(1'd0),
	.TXPRBSSEL(1'd0),
	.TXPRECURSOR(1'd0),
	.TXPRECURSORINV(1'd0),
	.TXRATE(1'd0),
	.TXRATEMODE(1'd0),
	.TXSEQUENCE(1'd0),
	.TXSTARTSEQ(1'd0),
	.TXSWING(1'd0),
	.TXSYNCALLIN(1'd0),
	.TXSYNCIN(1'd0),
	.TXSYNCMODE(1'd0),
	.TXSYSCLKSEL(1'd0),
	.TXUSERRDY(main_genericstandalone_tx_mmcm_locked),
	.TXUSRCLK(eth_tx_half_clk),
	.TXUSRCLK2(eth_tx_half_clk),
	.DRPDO(main_genericstandalone_drpdo),
	.DRPRDY(main_genericstandalone_drprdy),
	.GTPTXN(sfp_txn),
	.GTPTXP(sfp_txp),
	.RXCHARISK({main_genericstandalone_rx_data0[18], main_genericstandalone_rx_data0[8]}),
	.RXDATA({main_genericstandalone_rx_data0[17:10], main_genericstandalone_rx_data0[7:0]}),
	.RXDISPERR({main_genericstandalone_rx_data0[19], main_genericstandalone_rx_data0[9]}),
	.RXOUTCLK(main_genericstandalone_rxoutclk),
	.RXPMARESETDONE(main_genericstandalone_rx_pma_reset_done),
	.RXRESETDONE(main_genericstandalone_rx_reset_done),
	.TXOUTCLK(main_genericstandalone_txoutclk),
	.TXRESETDONE(main_genericstandalone_tx_reset_done)
);

BUFH BUFH_1(
	.I(main_genericstandalone_txoutclk),
	.O(main_genericstandalone_txoutclk_rebuffer)
);

BUFG BUFG_2(
	.I(main_genericstandalone_rxoutclk),
	.O(main_genericstandalone_rxoutclk_rebuffer)
);

MMCME2_BASE #(
	.CLKFBOUT_MULT_F(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE_F(5'd16),
	.CLKOUT1_DIVIDE(4'd8),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_BASE (
	.CLKFBIN(main_genericstandalone_tx_mmcm_fb),
	.CLKIN1(main_genericstandalone_txoutclk_rebuffer),
	.RST(main_genericstandalone_tx_mmcm_reset),
	.CLKFBOUT(main_genericstandalone_tx_mmcm_fb),
	.CLKOUT0(main_genericstandalone_clk_tx_half_unbuf),
	.CLKOUT1(main_genericstandalone_clk_tx_unbuf),
	.LOCKED(main_genericstandalone_tx_mmcm_locked)
);

BUFH BUFH_2(
	.I(main_genericstandalone_clk_tx_half_unbuf),
	.O(eth_tx_half_clk)
);

BUFH BUFH_3(
	.I(main_genericstandalone_clk_tx_unbuf),
	.O(eth_tx_clk)
);

MMCME2_BASE #(
	.CLKFBOUT_MULT_F(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE_F(5'd16),
	.CLKOUT1_DIVIDE(4'd8),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_BASE_1 (
	.CLKFBIN(main_genericstandalone_rx_mmcm_fb),
	.CLKIN1(main_genericstandalone_rxoutclk_rebuffer),
	.RST(main_genericstandalone_rx_mmcm_reset),
	.CLKFBOUT(main_genericstandalone_rx_mmcm_fb),
	.CLKOUT0(main_genericstandalone_clk_rx_half_unbuf),
	.CLKOUT1(main_genericstandalone_clk_rx_unbuf),
	.LOCKED(main_genericstandalone_rx_mmcm_locked)
);

BUFG BUFG_3(
	.I(main_genericstandalone_clk_rx_half_unbuf),
	.O(eth_rx_half_clk)
);

BUFG BUFG_4(
	.I(main_genericstandalone_clk_rx_unbuf),
	.O(eth_rx_clk)
);

reg [10:0] storage_2[0:4];
reg [10:0] memdat_2;
always @(posedge eth_rx_clk) begin : mem_write_block_7
	if (main_genericstandalone_crc32_checker_syncfifo_wrport_we)
		storage_2[main_genericstandalone_crc32_checker_syncfifo_wrport_adr] <= main_genericstandalone_crc32_checker_syncfifo_wrport_dat_w;
	memdat_2 <= storage_2[main_genericstandalone_crc32_checker_syncfifo_wrport_adr];
end

always @(posedge eth_rx_clk) begin : mem_write_block_8
end

assign main_genericstandalone_crc32_checker_syncfifo_wrport_dat_r = memdat_2;
assign main_genericstandalone_crc32_checker_syncfifo_rdport_dat_r = storage_2[main_genericstandalone_crc32_checker_syncfifo_rdport_adr];

reg [80:0] storage_3[0:63];
reg [5:0] memadr_3;
reg [5:0] memadr_4;
always @(posedge sys_clk) begin : mem_write_block_9
	if (main_genericstandalone_tx_cdc_wrport_we)
		storage_3[main_genericstandalone_tx_cdc_wrport_adr] <= main_genericstandalone_tx_cdc_wrport_dat_w;
	memadr_3 <= main_genericstandalone_tx_cdc_wrport_adr;
end

always @(posedge eth_tx_clk) begin : mem_write_block_10
	memadr_4 <= main_genericstandalone_tx_cdc_rdport_adr;
end

assign main_genericstandalone_tx_cdc_wrport_dat_r = storage_3[memadr_3];
assign main_genericstandalone_tx_cdc_rdport_dat_r = storage_3[memadr_4];

reg [80:0] storage_4[0:63];
reg [5:0] memadr_5;
reg [5:0] memadr_6;
always @(posedge eth_rx_clk) begin : mem_write_block_11
	if (main_genericstandalone_rx_cdc_wrport_we)
		storage_4[main_genericstandalone_rx_cdc_wrport_adr] <= main_genericstandalone_rx_cdc_wrport_dat_w;
	memadr_5 <= main_genericstandalone_rx_cdc_wrport_adr;
end

always @(posedge sys_clk) begin : mem_write_block_12
	memadr_6 <= main_genericstandalone_rx_cdc_rdport_adr;
end

assign main_genericstandalone_rx_cdc_wrport_dat_r = storage_4[memadr_5];
assign main_genericstandalone_rx_cdc_rdport_dat_r = storage_4[memadr_6];

reg [13:0] storage_5[0:3];
reg [13:0] memdat_3;
always @(posedge sys_clk) begin : mem_write_block_13
	if (main_genericstandalone_sram61_we)
		storage_5[main_genericstandalone_sram59_adr] <= main_genericstandalone_sram62_dat_w;
	memdat_3 <= storage_5[main_genericstandalone_sram59_adr];
end

always @(posedge sys_clk) begin : mem_write_block_14
end

assign main_genericstandalone_sram60_dat_r = memdat_3;
assign main_genericstandalone_sram65_dat_r = storage_5[main_genericstandalone_sram64_adr];

reg [63:0] mem_1[0:190];
reg [7:0] memadr_7;
reg [7:0] memadr_8;
always @(posedge sys_clk) begin : mem_write_block_15
	if (main_genericstandalone_sram74_we)
		mem_1[main_genericstandalone_sram72_adr] <= main_genericstandalone_sram75_dat_w;
	memadr_7 <= main_genericstandalone_sram72_adr;
end

always @(posedge sys_clk) begin : mem_write_block_16
	memadr_8 <= main_genericstandalone_sram0_adr;
end

assign main_genericstandalone_sram73_dat_r = mem_1[memadr_7];
assign main_genericstandalone_sram0_dat_r = mem_1[memadr_8];

reg [63:0] mem_2[0:190];
reg [7:0] memadr_9;
reg [7:0] memadr_10;
always @(posedge sys_clk) begin : mem_write_block_17
	if (main_genericstandalone_sram78_we)
		mem_2[main_genericstandalone_sram76_adr] <= main_genericstandalone_sram79_dat_w;
	memadr_9 <= main_genericstandalone_sram76_adr;
end

always @(posedge sys_clk) begin : mem_write_block_18
	memadr_10 <= main_genericstandalone_sram1_adr;
end

assign main_genericstandalone_sram77_dat_r = mem_2[memadr_9];
assign main_genericstandalone_sram1_dat_r = mem_2[memadr_10];

reg [63:0] mem_3[0:190];
reg [7:0] memadr_11;
reg [7:0] memadr_12;
always @(posedge sys_clk) begin : mem_write_block_19
	if (main_genericstandalone_sram82_we)
		mem_3[main_genericstandalone_sram80_adr] <= main_genericstandalone_sram83_dat_w;
	memadr_11 <= main_genericstandalone_sram80_adr;
end

always @(posedge sys_clk) begin : mem_write_block_20
	memadr_12 <= main_genericstandalone_sram2_adr;
end

assign main_genericstandalone_sram81_dat_r = mem_3[memadr_11];
assign main_genericstandalone_sram2_dat_r = mem_3[memadr_12];

reg [63:0] mem_4[0:190];
reg [7:0] memadr_13;
reg [7:0] memadr_14;
always @(posedge sys_clk) begin : mem_write_block_21
	if (main_genericstandalone_sram86_we)
		mem_4[main_genericstandalone_sram84_adr] <= main_genericstandalone_sram87_dat_w;
	memadr_13 <= main_genericstandalone_sram84_adr;
end

always @(posedge sys_clk) begin : mem_write_block_22
	memadr_14 <= main_genericstandalone_sram3_adr;
end

assign main_genericstandalone_sram85_dat_r = mem_4[memadr_13];
assign main_genericstandalone_sram3_dat_r = mem_4[memadr_14];

reg [13:0] storage_6[0:3];
reg [13:0] memdat_4;
always @(posedge sys_clk) begin : mem_write_block_23
	if (main_genericstandalone_sram141_we)
		storage_6[main_genericstandalone_sram139_adr] <= main_genericstandalone_sram142_dat_w;
	memdat_4 <= storage_6[main_genericstandalone_sram139_adr];
end

always @(posedge sys_clk) begin : mem_write_block_24
end

assign main_genericstandalone_sram140_dat_r = memdat_4;
assign main_genericstandalone_sram145_dat_r = storage_6[main_genericstandalone_sram144_adr];

VexRiscv_G VexRiscv_G(
	.clk(sys_kernel_clk),
	.dBusWishbone_ACK(main_genericstandalone_kernel_cpu_dbus_ack),
	.dBusWishbone_DAT_MISO(main_genericstandalone_kernel_cpu_dbus_dat_r),
	.dBusWishbone_ERR(main_genericstandalone_kernel_cpu_dbus_err),
	.externalInterruptArray(main_genericstandalone_kernel_cpu_interrupt),
	.externalResetVector(31'd1157627904),
	.iBusWishbone_ACK(main_genericstandalone_kernel_cpu_ibus_ack),
	.iBusWishbone_DAT_MISO(main_genericstandalone_kernel_cpu_ibus_dat_r),
	.iBusWishbone_ERR(main_genericstandalone_kernel_cpu_ibus_err),
	.reset(sys_kernel_rst),
	.timerInterrupt(1'd0),
	.dBusWishbone_ADR(main_genericstandalone_kernel_cpu_dbus_adr),
	.dBusWishbone_BTE(main_genericstandalone_kernel_cpu_dbus_bte),
	.dBusWishbone_CTI(main_genericstandalone_kernel_cpu_dbus_cti),
	.dBusWishbone_CYC(main_genericstandalone_kernel_cpu_dbus_cyc),
	.dBusWishbone_DAT_MOSI(main_genericstandalone_kernel_cpu_dbus_dat_w),
	.dBusWishbone_SEL(main_genericstandalone_kernel_cpu_dbus_sel),
	.dBusWishbone_STB(main_genericstandalone_kernel_cpu_dbus_stb),
	.dBusWishbone_WE(main_genericstandalone_kernel_cpu_dbus_we),
	.iBusWishbone_ADR(main_genericstandalone_kernel_cpu_ibus_adr),
	.iBusWishbone_BTE(main_genericstandalone_kernel_cpu_ibus_bte),
	.iBusWishbone_CTI(main_genericstandalone_kernel_cpu_ibus_cti),
	.iBusWishbone_CYC(main_genericstandalone_kernel_cpu_ibus_cyc),
	.iBusWishbone_DAT_MOSI(main_genericstandalone_kernel_cpu_ibus_dat_w),
	.iBusWishbone_SEL(main_genericstandalone_kernel_cpu_ibus_sel),
	.iBusWishbone_STB(main_genericstandalone_kernel_cpu_ibus_stb),
	.iBusWishbone_WE(main_genericstandalone_kernel_cpu_ibus_we)
);

ROM256X1 #(
	.INIT(24'd10176178)
) identifier_str0 (
	.A0(main_genericstandalone_add_identifier_storage[0]),
	.A1(main_genericstandalone_add_identifier_storage[1]),
	.A2(main_genericstandalone_add_identifier_storage[2]),
	.A3(main_genericstandalone_add_identifier_storage[3]),
	.A4(main_genericstandalone_add_identifier_storage[4]),
	.A5(main_genericstandalone_add_identifier_storage[5]),
	.A6(main_genericstandalone_add_identifier_storage[6]),
	.A7(main_genericstandalone_add_identifier_storage[7]),
	.O(main_genericstandalone_add_identifier_status[0])
);

ROM256X1 #(
	.INIT(23'd5390292)
) identifier_str1 (
	.A0(main_genericstandalone_add_identifier_storage[0]),
	.A1(main_genericstandalone_add_identifier_storage[1]),
	.A2(main_genericstandalone_add_identifier_storage[2]),
	.A3(main_genericstandalone_add_identifier_storage[3]),
	.A4(main_genericstandalone_add_identifier_storage[4]),
	.A5(main_genericstandalone_add_identifier_storage[5]),
	.A6(main_genericstandalone_add_identifier_storage[6]),
	.A7(main_genericstandalone_add_identifier_storage[7]),
	.O(main_genericstandalone_add_identifier_status[1])
);

ROM256X1 #(
	.INIT(25'd28106596)
) identifier_str2 (
	.A0(main_genericstandalone_add_identifier_storage[0]),
	.A1(main_genericstandalone_add_identifier_storage[1]),
	.A2(main_genericstandalone_add_identifier_storage[2]),
	.A3(main_genericstandalone_add_identifier_storage[3]),
	.A4(main_genericstandalone_add_identifier_storage[4]),
	.A5(main_genericstandalone_add_identifier_storage[5]),
	.A6(main_genericstandalone_add_identifier_storage[6]),
	.A7(main_genericstandalone_add_identifier_storage[7]),
	.O(main_genericstandalone_add_identifier_status[2])
);

ROM256X1 #(
	.INIT(18'd138199)
) identifier_str3 (
	.A0(main_genericstandalone_add_identifier_storage[0]),
	.A1(main_genericstandalone_add_identifier_storage[1]),
	.A2(main_genericstandalone_add_identifier_storage[2]),
	.A3(main_genericstandalone_add_identifier_storage[3]),
	.A4(main_genericstandalone_add_identifier_storage[4]),
	.A5(main_genericstandalone_add_identifier_storage[5]),
	.A6(main_genericstandalone_add_identifier_storage[6]),
	.A7(main_genericstandalone_add_identifier_storage[7]),
	.O(main_genericstandalone_add_identifier_status[3])
);

ROM256X1 #(
	.INIT(22'd3572779)
) identifier_str4 (
	.A0(main_genericstandalone_add_identifier_storage[0]),
	.A1(main_genericstandalone_add_identifier_storage[1]),
	.A2(main_genericstandalone_add_identifier_storage[2]),
	.A3(main_genericstandalone_add_identifier_storage[3]),
	.A4(main_genericstandalone_add_identifier_storage[4]),
	.A5(main_genericstandalone_add_identifier_storage[5]),
	.A6(main_genericstandalone_add_identifier_storage[6]),
	.A7(main_genericstandalone_add_identifier_storage[7]),
	.O(main_genericstandalone_add_identifier_status[4])
);

ROM256X1 #(
	.INIT(25'd33554430)
) identifier_str5 (
	.A0(main_genericstandalone_add_identifier_storage[0]),
	.A1(main_genericstandalone_add_identifier_storage[1]),
	.A2(main_genericstandalone_add_identifier_storage[2]),
	.A3(main_genericstandalone_add_identifier_storage[3]),
	.A4(main_genericstandalone_add_identifier_storage[4]),
	.A5(main_genericstandalone_add_identifier_storage[5]),
	.A6(main_genericstandalone_add_identifier_storage[6]),
	.A7(main_genericstandalone_add_identifier_storage[7]),
	.O(main_genericstandalone_add_identifier_status[5])
);

ROM256X1 #(
	.INIT(25'd33419232)
) identifier_str6 (
	.A0(main_genericstandalone_add_identifier_storage[0]),
	.A1(main_genericstandalone_add_identifier_storage[1]),
	.A2(main_genericstandalone_add_identifier_storage[2]),
	.A3(main_genericstandalone_add_identifier_storage[3]),
	.A4(main_genericstandalone_add_identifier_storage[4]),
	.A5(main_genericstandalone_add_identifier_storage[5]),
	.A6(main_genericstandalone_add_identifier_storage[6]),
	.A7(main_genericstandalone_add_identifier_storage[7]),
	.O(main_genericstandalone_add_identifier_status[6])
);

ROM256X1 #(
	.INIT(1'd0)
) identifier_str7 (
	.A0(main_genericstandalone_add_identifier_storage[0]),
	.A1(main_genericstandalone_add_identifier_storage[1]),
	.A2(main_genericstandalone_add_identifier_storage[2]),
	.A3(main_genericstandalone_add_identifier_storage[3]),
	.A4(main_genericstandalone_add_identifier_storage[4]),
	.A5(main_genericstandalone_add_identifier_storage[5]),
	.A6(main_genericstandalone_add_identifier_storage[6]),
	.A7(main_genericstandalone_add_identifier_storage[7]),
	.O(main_genericstandalone_add_identifier_status[7])
);

IBUFDS_GTE2 #(
	.CLKCM_CFG("TRUE"),
	.CLKRCV_TRST("TRUE"),
	.CLKSWING_CFG(2'd3)
) IBUFDS_GTE2_1 (
	.CEB(1'd0),
	.I(cdr_clk_clean_p),
	.IB(cdr_clk_clean_n),
	.O(main_genericstandalone_cdr_clk)
);

BUFG BUFG_5(
	.I(main_genericstandalone_cdr_clk),
	.O(main_genericstandalone_cdr_clk_buf)
);

MMCME2_ADV #(
	.CLKFBOUT_MULT_F(4'd8),
	.CLKIN1_PERIOD(8.0),
	.CLKIN2_PERIOD(8.0),
	.CLKOUT0_DIVIDE_F(4'd8),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(2'd2),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(2'd2),
	.CLKOUT2_PHASE(90.0),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_ADV (
	.CLKFBIN(main_genericstandalone_rtiosyscrg_mmcm_fb_in),
	.CLKIN1(main_genericstandalone_cdr_clk_buf),
	.CLKIN2(bootstrap_clk),
	.CLKINSEL(main_genericstandalone_genericstandalone_crg_o_clk_sw),
	.RST(main_genericstandalone_genericstandalone_crg_o_reset),
	.CLKFBOUT(main_genericstandalone_rtiosyscrg_mmcm_fb_out),
	.CLKOUT0(main_genericstandalone_rtiosyscrg_mmcm_sys),
	.CLKOUT1(main_genericstandalone_rtiosyscrg_mmcm_sys4x),
	.CLKOUT2(main_genericstandalone_rtiosyscrg_mmcm_sys4x_dqs),
	.LOCKED(main_genericstandalone_rtiosyscrg_mmcm_locked)
);

BUFG BUFG_6(
	.I(main_genericstandalone_rtiosyscrg_mmcm_sys),
	.O(sys_clk)
);

BUFG BUFG_7(
	.I(main_genericstandalone_rtiosyscrg_mmcm_sys4x),
	.O(sys4x_clk)
);

BUFG BUFG_8(
	.I(main_genericstandalone_rtiosyscrg_mmcm_fb_out),
	.O(main_genericstandalone_rtiosyscrg_mmcm_fb_in)
);

BUFG BUFG_9(
	.I(main_genericstandalone_rtiosyscrg_mmcm_sys4x_dqs),
	.O(sys4x_dqs_clk)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(main_genericstandalone_rtiosyscrg_async_reset),
	.Q(main_genericstandalone_rtiosyscrg_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(sys_clk),
	.CE(1'd1),
	.D(main_genericstandalone_rtiosyscrg_rst_meta),
	.PRE(main_genericstandalone_rtiosyscrg_async_reset),
	.Q(main_genericstandalone_rtiosyscrg_rst_unbuf)
);

BUFG BUFG_10(
	.I(main_genericstandalone_rtiosyscrg_rst_unbuf),
	.O(sys_rst)
);

IBUFDS IBUFDS(
	.I(sma_clkin_p),
	.IB(sma_clkin_n),
	.O(main_genericstandalone_sma_clkin_se)
);

BUFIO BUFIO(
	.I(main_genericstandalone_sma_clkin_se),
	.O(main_genericstandalone_sma_clkin_buffered)
);

ODDR ODDR(
	.C(main_genericstandalone_sma_clkin_buffered),
	.CE(1'd1),
	.D1(1'd0),
	.D2(1'd1),
	.Q(main_genericstandalone_cdr_clk_se)
);

OBUFDS OBUFDS_1(
	.I(main_genericstandalone_cdr_clk_se),
	.O(cdr_clk_p),
	.OB(cdr_clk_n)
);

assign i2c_scl = main_genericstandalone_i2c_tstriple0_oe ? main_genericstandalone_i2c_tstriple0_o : 1'bz;
assign main_genericstandalone_i2c_tstriple0_i = i2c_scl;

assign i2c_sda = main_genericstandalone_i2c_tstriple1_oe ? main_genericstandalone_i2c_tstriple1_o : 1'bz;
assign main_genericstandalone_i2c_tstriple1_i = i2c_sda;

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_16 (
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x0_serdes_ser_in),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x0_serdes_i1[7]),
	.Q2(main_inout_8x0_serdes_i1[6]),
	.Q3(main_inout_8x0_serdes_i1[5]),
	.Q4(main_inout_8x0_serdes_i1[4]),
	.Q5(main_inout_8x0_serdes_i1[3]),
	.Q6(main_inout_8x0_serdes_i1[2]),
	.Q7(main_inout_8x0_serdes_i1[1]),
	.Q8(main_inout_8x0_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_45 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x0_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x0_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x0_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x0_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x0_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x0_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x0_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x0_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x0_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x0_serdes_ser_out),
	.TQ(main_inout_8x0_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE (
	.I(main_inout_8x0_serdes_ser_out),
	.IBUFDISABLE((~main_inout_8x0_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x0_serdes_t_out)),
	.T(main_inout_8x0_serdes_t_out),
	.IO(dio0_p),
	.IOB(dio0_n),
	.O(main_inout_8x0_serdes_ser_in)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_17 (
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x1_serdes_ser_in),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x1_serdes_i1[7]),
	.Q2(main_inout_8x1_serdes_i1[6]),
	.Q3(main_inout_8x1_serdes_i1[5]),
	.Q4(main_inout_8x1_serdes_i1[4]),
	.Q5(main_inout_8x1_serdes_i1[3]),
	.Q6(main_inout_8x1_serdes_i1[2]),
	.Q7(main_inout_8x1_serdes_i1[1]),
	.Q8(main_inout_8x1_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_46 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x1_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x1_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x1_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x1_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x1_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x1_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x1_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x1_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x1_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x1_serdes_ser_out),
	.TQ(main_inout_8x1_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_1 (
	.I(main_inout_8x1_serdes_ser_out),
	.IBUFDISABLE((~main_inout_8x1_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x1_serdes_t_out)),
	.T(main_inout_8x1_serdes_t_out),
	.IO(dio0_p_1),
	.IOB(dio0_n_1),
	.O(main_inout_8x1_serdes_ser_in)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_18 (
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x2_serdes_ser_in),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x2_serdes_i1[7]),
	.Q2(main_inout_8x2_serdes_i1[6]),
	.Q3(main_inout_8x2_serdes_i1[5]),
	.Q4(main_inout_8x2_serdes_i1[4]),
	.Q5(main_inout_8x2_serdes_i1[3]),
	.Q6(main_inout_8x2_serdes_i1[2]),
	.Q7(main_inout_8x2_serdes_i1[1]),
	.Q8(main_inout_8x2_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_47 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x2_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x2_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x2_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x2_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x2_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x2_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x2_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x2_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x2_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x2_serdes_ser_out),
	.TQ(main_inout_8x2_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_2 (
	.I(main_inout_8x2_serdes_ser_out),
	.IBUFDISABLE((~main_inout_8x2_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x2_serdes_t_out)),
	.T(main_inout_8x2_serdes_t_out),
	.IO(dio0_p_2),
	.IOB(dio0_n_2),
	.O(main_inout_8x2_serdes_ser_in)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_19 (
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x3_serdes_ser_in),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x3_serdes_i1[7]),
	.Q2(main_inout_8x3_serdes_i1[6]),
	.Q3(main_inout_8x3_serdes_i1[5]),
	.Q4(main_inout_8x3_serdes_i1[4]),
	.Q5(main_inout_8x3_serdes_i1[3]),
	.Q6(main_inout_8x3_serdes_i1[2]),
	.Q7(main_inout_8x3_serdes_i1[1]),
	.Q8(main_inout_8x3_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_48 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x3_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x3_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x3_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x3_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x3_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x3_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x3_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x3_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x3_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x3_serdes_ser_out),
	.TQ(main_inout_8x3_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_3 (
	.I(main_inout_8x3_serdes_ser_out),
	.IBUFDISABLE((~main_inout_8x3_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x3_serdes_t_out)),
	.T(main_inout_8x3_serdes_t_out),
	.IO(dio0_p_3),
	.IOB(dio0_n_3),
	.O(main_inout_8x3_serdes_ser_in)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_49 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x0_o0[0] ^ 1'd0)),
	.D2((main_output_8x0_o0[1] ^ 1'd0)),
	.D3((main_output_8x0_o0[2] ^ 1'd0)),
	.D4((main_output_8x0_o0[3] ^ 1'd0)),
	.D5((main_output_8x0_o0[4] ^ 1'd0)),
	.D6((main_output_8x0_o0[5] ^ 1'd0)),
	.D7((main_output_8x0_o0[6] ^ 1'd0)),
	.D8((main_output_8x0_o0[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x0_t_in0),
	.TCE(1'd1),
	.OQ(main_output_8x0_ser_out0),
	.TQ(main_output_8x0_t_out0)
);

IOBUFDS IOBUFDS(
	.I(main_output_8x0_ser_out0),
	.T(main_output_8x0_t_out0),
	.IO(dio0_p_4),
	.IOB(dio0_n_4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_50 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x1_o0[0] ^ 1'd0)),
	.D2((main_output_8x1_o0[1] ^ 1'd0)),
	.D3((main_output_8x1_o0[2] ^ 1'd0)),
	.D4((main_output_8x1_o0[3] ^ 1'd0)),
	.D5((main_output_8x1_o0[4] ^ 1'd0)),
	.D6((main_output_8x1_o0[5] ^ 1'd0)),
	.D7((main_output_8x1_o0[6] ^ 1'd0)),
	.D8((main_output_8x1_o0[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x1_t_in0),
	.TCE(1'd1),
	.OQ(main_output_8x1_ser_out0),
	.TQ(main_output_8x1_t_out0)
);

IOBUFDS IOBUFDS_1(
	.I(main_output_8x1_ser_out0),
	.T(main_output_8x1_t_out0),
	.IO(dio0_p_5),
	.IOB(dio0_n_5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_51 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x2_o[0] ^ 1'd0)),
	.D2((main_output_8x2_o[1] ^ 1'd0)),
	.D3((main_output_8x2_o[2] ^ 1'd0)),
	.D4((main_output_8x2_o[3] ^ 1'd0)),
	.D5((main_output_8x2_o[4] ^ 1'd0)),
	.D6((main_output_8x2_o[5] ^ 1'd0)),
	.D7((main_output_8x2_o[6] ^ 1'd0)),
	.D8((main_output_8x2_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x2_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x2_ser_out),
	.TQ(main_output_8x2_t_out)
);

IOBUFDS IOBUFDS_2(
	.I(main_output_8x2_ser_out),
	.T(main_output_8x2_t_out),
	.IO(dio0_p_6),
	.IOB(dio0_n_6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_52 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x3_o[0] ^ 1'd0)),
	.D2((main_output_8x3_o[1] ^ 1'd0)),
	.D3((main_output_8x3_o[2] ^ 1'd0)),
	.D4((main_output_8x3_o[3] ^ 1'd0)),
	.D5((main_output_8x3_o[4] ^ 1'd0)),
	.D6((main_output_8x3_o[5] ^ 1'd0)),
	.D7((main_output_8x3_o[6] ^ 1'd0)),
	.D8((main_output_8x3_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x3_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x3_ser_out),
	.TQ(main_output_8x3_t_out)
);

IOBUFDS IOBUFDS_3(
	.I(main_output_8x3_ser_out),
	.T(main_output_8x3_t_out),
	.IO(dio0_p_7),
	.IOB(dio0_n_7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_53 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x4_o[0] ^ 1'd0)),
	.D2((main_output_8x4_o[1] ^ 1'd0)),
	.D3((main_output_8x4_o[2] ^ 1'd0)),
	.D4((main_output_8x4_o[3] ^ 1'd0)),
	.D5((main_output_8x4_o[4] ^ 1'd0)),
	.D6((main_output_8x4_o[5] ^ 1'd0)),
	.D7((main_output_8x4_o[6] ^ 1'd0)),
	.D8((main_output_8x4_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x4_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x4_ser_out),
	.TQ(main_output_8x4_t_out)
);

IOBUFDS IOBUFDS_4(
	.I(main_output_8x4_ser_out),
	.T(main_output_8x4_t_out),
	.IO(dio1_p),
	.IOB(dio1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_54 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x5_o[0] ^ 1'd0)),
	.D2((main_output_8x5_o[1] ^ 1'd0)),
	.D3((main_output_8x5_o[2] ^ 1'd0)),
	.D4((main_output_8x5_o[3] ^ 1'd0)),
	.D5((main_output_8x5_o[4] ^ 1'd0)),
	.D6((main_output_8x5_o[5] ^ 1'd0)),
	.D7((main_output_8x5_o[6] ^ 1'd0)),
	.D8((main_output_8x5_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x5_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x5_ser_out),
	.TQ(main_output_8x5_t_out)
);

IOBUFDS IOBUFDS_5(
	.I(main_output_8x5_ser_out),
	.T(main_output_8x5_t_out),
	.IO(dio1_p_1),
	.IOB(dio1_n_1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_55 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x6_o[0] ^ 1'd0)),
	.D2((main_output_8x6_o[1] ^ 1'd0)),
	.D3((main_output_8x6_o[2] ^ 1'd0)),
	.D4((main_output_8x6_o[3] ^ 1'd0)),
	.D5((main_output_8x6_o[4] ^ 1'd0)),
	.D6((main_output_8x6_o[5] ^ 1'd0)),
	.D7((main_output_8x6_o[6] ^ 1'd0)),
	.D8((main_output_8x6_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x6_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x6_ser_out),
	.TQ(main_output_8x6_t_out)
);

IOBUFDS IOBUFDS_6(
	.I(main_output_8x6_ser_out),
	.T(main_output_8x6_t_out),
	.IO(dio1_p_2),
	.IOB(dio1_n_2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_56 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x7_o[0] ^ 1'd0)),
	.D2((main_output_8x7_o[1] ^ 1'd0)),
	.D3((main_output_8x7_o[2] ^ 1'd0)),
	.D4((main_output_8x7_o[3] ^ 1'd0)),
	.D5((main_output_8x7_o[4] ^ 1'd0)),
	.D6((main_output_8x7_o[5] ^ 1'd0)),
	.D7((main_output_8x7_o[6] ^ 1'd0)),
	.D8((main_output_8x7_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x7_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x7_ser_out),
	.TQ(main_output_8x7_t_out)
);

IOBUFDS IOBUFDS_7(
	.I(main_output_8x7_ser_out),
	.T(main_output_8x7_t_out),
	.IO(dio1_p_3),
	.IOB(dio1_n_3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_57 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x8_o[0] ^ 1'd0)),
	.D2((main_output_8x8_o[1] ^ 1'd0)),
	.D3((main_output_8x8_o[2] ^ 1'd0)),
	.D4((main_output_8x8_o[3] ^ 1'd0)),
	.D5((main_output_8x8_o[4] ^ 1'd0)),
	.D6((main_output_8x8_o[5] ^ 1'd0)),
	.D7((main_output_8x8_o[6] ^ 1'd0)),
	.D8((main_output_8x8_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x8_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x8_ser_out),
	.TQ(main_output_8x8_t_out)
);

IOBUFDS IOBUFDS_8(
	.I(main_output_8x8_ser_out),
	.T(main_output_8x8_t_out),
	.IO(dio1_p_4),
	.IOB(dio1_n_4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_58 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x9_o[0] ^ 1'd0)),
	.D2((main_output_8x9_o[1] ^ 1'd0)),
	.D3((main_output_8x9_o[2] ^ 1'd0)),
	.D4((main_output_8x9_o[3] ^ 1'd0)),
	.D5((main_output_8x9_o[4] ^ 1'd0)),
	.D6((main_output_8x9_o[5] ^ 1'd0)),
	.D7((main_output_8x9_o[6] ^ 1'd0)),
	.D8((main_output_8x9_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x9_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x9_ser_out),
	.TQ(main_output_8x9_t_out)
);

IOBUFDS IOBUFDS_9(
	.I(main_output_8x9_ser_out),
	.T(main_output_8x9_t_out),
	.IO(dio1_p_5),
	.IOB(dio1_n_5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_59 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x10_o[0] ^ 1'd0)),
	.D2((main_output_8x10_o[1] ^ 1'd0)),
	.D3((main_output_8x10_o[2] ^ 1'd0)),
	.D4((main_output_8x10_o[3] ^ 1'd0)),
	.D5((main_output_8x10_o[4] ^ 1'd0)),
	.D6((main_output_8x10_o[5] ^ 1'd0)),
	.D7((main_output_8x10_o[6] ^ 1'd0)),
	.D8((main_output_8x10_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x10_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x10_ser_out),
	.TQ(main_output_8x10_t_out)
);

IOBUFDS IOBUFDS_10(
	.I(main_output_8x10_ser_out),
	.T(main_output_8x10_t_out),
	.IO(dio1_p_6),
	.IOB(dio1_n_6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_60 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x11_o[0] ^ 1'd0)),
	.D2((main_output_8x11_o[1] ^ 1'd0)),
	.D3((main_output_8x11_o[2] ^ 1'd0)),
	.D4((main_output_8x11_o[3] ^ 1'd0)),
	.D5((main_output_8x11_o[4] ^ 1'd0)),
	.D6((main_output_8x11_o[5] ^ 1'd0)),
	.D7((main_output_8x11_o[6] ^ 1'd0)),
	.D8((main_output_8x11_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x11_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x11_ser_out),
	.TQ(main_output_8x11_t_out)
);

IOBUFDS IOBUFDS_11(
	.I(main_output_8x11_ser_out),
	.T(main_output_8x11_t_out),
	.IO(dio1_p_7),
	.IOB(dio1_n_7)
);

OBUFTDS OBUFTDS_2(
	.I(main_spimaster0_interface_cs1[0]),
	.T(main_spimaster0_interface_offline0),
	.O(urukul2_spi_p_cs_n[0]),
	.OB(urukul2_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_3(
	.I(main_spimaster0_interface_cs1[1]),
	.T(main_spimaster0_interface_offline0),
	.O(urukul2_spi_p_cs_n[1]),
	.OB(urukul2_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_4(
	.I(main_spimaster0_interface_cs1[2]),
	.T(main_spimaster0_interface_offline0),
	.O(urukul2_spi_p_cs_n[2]),
	.OB(urukul2_spi_n_cs_n[2])
);

OBUFTDS OBUFTDS_5(
	.I(main_spimaster0_interface_clk0),
	.T(main_spimaster0_interface_offline0),
	.O(urukul2_spi_p_clk),
	.OB(urukul2_spi_n_clk)
);

IOBUFDS IOBUFDS_12(
	.I(main_spimaster0_interface_sdo0),
	.T((main_spimaster0_interface_offline0 | main_spimaster0_interface_half_duplex0)),
	.IO(urukul2_spi_p_mosi),
	.IOB(urukul2_spi_n_mosi),
	.O(main_spimaster0_interface_mosi0)
);

IOBUFDS IOBUFDS_13(
	.I(main_spimaster0_interface_sdo0),
	.T(1'd1),
	.IO(urukul2_spi_p_miso),
	.IOB(urukul2_spi_n_miso),
	.O(main_spimaster0_interface_miso0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_61 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x0_o1[0] ^ 1'd0)),
	.D2((main_output_8x0_o1[1] ^ 1'd0)),
	.D3((main_output_8x0_o1[2] ^ 1'd0)),
	.D4((main_output_8x0_o1[3] ^ 1'd0)),
	.D5((main_output_8x0_o1[4] ^ 1'd0)),
	.D6((main_output_8x0_o1[5] ^ 1'd0)),
	.D7((main_output_8x0_o1[6] ^ 1'd0)),
	.D8((main_output_8x0_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x0_t_in1),
	.TCE(1'd1),
	.OQ(main_output_8x0_ser_out1),
	.TQ(main_output_8x0_t_out1)
);

IOBUFDS IOBUFDS_14(
	.I(main_output_8x0_ser_out1),
	.T(main_output_8x0_t_out1),
	.IO(urukul2_io_update_p),
	.IOB(urukul2_io_update_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_62 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x12_o[0] ^ 1'd0)),
	.D2((main_output_8x12_o[1] ^ 1'd0)),
	.D3((main_output_8x12_o[2] ^ 1'd0)),
	.D4((main_output_8x12_o[3] ^ 1'd0)),
	.D5((main_output_8x12_o[4] ^ 1'd0)),
	.D6((main_output_8x12_o[5] ^ 1'd0)),
	.D7((main_output_8x12_o[6] ^ 1'd0)),
	.D8((main_output_8x12_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x12_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x12_ser_out),
	.TQ(main_output_8x12_t_out)
);

IOBUFDS IOBUFDS_15(
	.I(main_output_8x12_ser_out),
	.T(main_output_8x12_t_out),
	.IO(urukul2_sw0_p),
	.IOB(urukul2_sw0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_63 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x13_o[0] ^ 1'd0)),
	.D2((main_output_8x13_o[1] ^ 1'd0)),
	.D3((main_output_8x13_o[2] ^ 1'd0)),
	.D4((main_output_8x13_o[3] ^ 1'd0)),
	.D5((main_output_8x13_o[4] ^ 1'd0)),
	.D6((main_output_8x13_o[5] ^ 1'd0)),
	.D7((main_output_8x13_o[6] ^ 1'd0)),
	.D8((main_output_8x13_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x13_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x13_ser_out),
	.TQ(main_output_8x13_t_out)
);

IOBUFDS IOBUFDS_16(
	.I(main_output_8x13_ser_out),
	.T(main_output_8x13_t_out),
	.IO(urukul2_sw1_p),
	.IOB(urukul2_sw1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_64 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x14_o[0] ^ 1'd0)),
	.D2((main_output_8x14_o[1] ^ 1'd0)),
	.D3((main_output_8x14_o[2] ^ 1'd0)),
	.D4((main_output_8x14_o[3] ^ 1'd0)),
	.D5((main_output_8x14_o[4] ^ 1'd0)),
	.D6((main_output_8x14_o[5] ^ 1'd0)),
	.D7((main_output_8x14_o[6] ^ 1'd0)),
	.D8((main_output_8x14_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x14_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x14_ser_out),
	.TQ(main_output_8x14_t_out)
);

IOBUFDS IOBUFDS_17(
	.I(main_output_8x14_ser_out),
	.T(main_output_8x14_t_out),
	.IO(urukul2_sw2_p),
	.IOB(urukul2_sw2_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_65 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x15_o[0] ^ 1'd0)),
	.D2((main_output_8x15_o[1] ^ 1'd0)),
	.D3((main_output_8x15_o[2] ^ 1'd0)),
	.D4((main_output_8x15_o[3] ^ 1'd0)),
	.D5((main_output_8x15_o[4] ^ 1'd0)),
	.D6((main_output_8x15_o[5] ^ 1'd0)),
	.D7((main_output_8x15_o[6] ^ 1'd0)),
	.D8((main_output_8x15_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x15_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x15_ser_out),
	.TQ(main_output_8x15_t_out)
);

IOBUFDS IOBUFDS_18(
	.I(main_output_8x15_ser_out),
	.T(main_output_8x15_t_out),
	.IO(urukul2_sw3_p),
	.IOB(urukul2_sw3_n)
);

OBUFTDS OBUFTDS_6(
	.I(main_spimaster1_interface_cs1[0]),
	.T(main_spimaster1_interface_offline0),
	.O(urukul4_spi_p_cs_n[0]),
	.OB(urukul4_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_7(
	.I(main_spimaster1_interface_cs1[1]),
	.T(main_spimaster1_interface_offline0),
	.O(urukul4_spi_p_cs_n[1]),
	.OB(urukul4_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_8(
	.I(main_spimaster1_interface_cs1[2]),
	.T(main_spimaster1_interface_offline0),
	.O(urukul4_spi_p_cs_n[2]),
	.OB(urukul4_spi_n_cs_n[2])
);

OBUFTDS OBUFTDS_9(
	.I(main_spimaster1_interface_clk0),
	.T(main_spimaster1_interface_offline0),
	.O(urukul4_spi_p_clk),
	.OB(urukul4_spi_n_clk)
);

IOBUFDS IOBUFDS_19(
	.I(main_spimaster1_interface_sdo0),
	.T((main_spimaster1_interface_offline0 | main_spimaster1_interface_half_duplex0)),
	.IO(urukul4_spi_p_mosi),
	.IOB(urukul4_spi_n_mosi),
	.O(main_spimaster1_interface_mosi0)
);

IOBUFDS IOBUFDS_20(
	.I(main_spimaster1_interface_sdo0),
	.T(1'd1),
	.IO(urukul4_spi_p_miso),
	.IOB(urukul4_spi_n_miso),
	.O(main_spimaster1_interface_miso0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_66 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x1_o1[0] ^ 1'd0)),
	.D2((main_output_8x1_o1[1] ^ 1'd0)),
	.D3((main_output_8x1_o1[2] ^ 1'd0)),
	.D4((main_output_8x1_o1[3] ^ 1'd0)),
	.D5((main_output_8x1_o1[4] ^ 1'd0)),
	.D6((main_output_8x1_o1[5] ^ 1'd0)),
	.D7((main_output_8x1_o1[6] ^ 1'd0)),
	.D8((main_output_8x1_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x1_t_in1),
	.TCE(1'd1),
	.OQ(main_output_8x1_ser_out1),
	.TQ(main_output_8x1_t_out1)
);

IOBUFDS IOBUFDS_21(
	.I(main_output_8x1_ser_out1),
	.T(main_output_8x1_t_out1),
	.IO(urukul4_io_update_p),
	.IOB(urukul4_io_update_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_67 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x16_o[0] ^ 1'd0)),
	.D2((main_output_8x16_o[1] ^ 1'd0)),
	.D3((main_output_8x16_o[2] ^ 1'd0)),
	.D4((main_output_8x16_o[3] ^ 1'd0)),
	.D5((main_output_8x16_o[4] ^ 1'd0)),
	.D6((main_output_8x16_o[5] ^ 1'd0)),
	.D7((main_output_8x16_o[6] ^ 1'd0)),
	.D8((main_output_8x16_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x16_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x16_ser_out),
	.TQ(main_output_8x16_t_out)
);

IOBUFDS IOBUFDS_22(
	.I(main_output_8x16_ser_out),
	.T(main_output_8x16_t_out),
	.IO(urukul4_sw0_p),
	.IOB(urukul4_sw0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_68 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x17_o[0] ^ 1'd0)),
	.D2((main_output_8x17_o[1] ^ 1'd0)),
	.D3((main_output_8x17_o[2] ^ 1'd0)),
	.D4((main_output_8x17_o[3] ^ 1'd0)),
	.D5((main_output_8x17_o[4] ^ 1'd0)),
	.D6((main_output_8x17_o[5] ^ 1'd0)),
	.D7((main_output_8x17_o[6] ^ 1'd0)),
	.D8((main_output_8x17_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x17_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x17_ser_out),
	.TQ(main_output_8x17_t_out)
);

IOBUFDS IOBUFDS_23(
	.I(main_output_8x17_ser_out),
	.T(main_output_8x17_t_out),
	.IO(urukul4_sw1_p),
	.IOB(urukul4_sw1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_69 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x18_o[0] ^ 1'd0)),
	.D2((main_output_8x18_o[1] ^ 1'd0)),
	.D3((main_output_8x18_o[2] ^ 1'd0)),
	.D4((main_output_8x18_o[3] ^ 1'd0)),
	.D5((main_output_8x18_o[4] ^ 1'd0)),
	.D6((main_output_8x18_o[5] ^ 1'd0)),
	.D7((main_output_8x18_o[6] ^ 1'd0)),
	.D8((main_output_8x18_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x18_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x18_ser_out),
	.TQ(main_output_8x18_t_out)
);

IOBUFDS IOBUFDS_24(
	.I(main_output_8x18_ser_out),
	.T(main_output_8x18_t_out),
	.IO(urukul4_sw2_p),
	.IOB(urukul4_sw2_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_70 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x19_o[0] ^ 1'd0)),
	.D2((main_output_8x19_o[1] ^ 1'd0)),
	.D3((main_output_8x19_o[2] ^ 1'd0)),
	.D4((main_output_8x19_o[3] ^ 1'd0)),
	.D5((main_output_8x19_o[4] ^ 1'd0)),
	.D6((main_output_8x19_o[5] ^ 1'd0)),
	.D7((main_output_8x19_o[6] ^ 1'd0)),
	.D8((main_output_8x19_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x19_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x19_ser_out),
	.TQ(main_output_8x19_t_out)
);

IOBUFDS IOBUFDS_25(
	.I(main_output_8x19_ser_out),
	.T(main_output_8x19_t_out),
	.IO(urukul4_sw3_p),
	.IOB(urukul4_sw3_n)
);

OBUFTDS OBUFTDS_10(
	.I(main_spimaster0_interface_clk1),
	.T(main_spimaster0_interface_offline1),
	.O(sampler6_adc_spi_p_clk),
	.OB(sampler6_adc_spi_n_clk)
);

IOBUFDS IOBUFDS_26(
	.I(main_spimaster0_interface_sdo1),
	.T(1'd1),
	.IO(sampler6_adc_spi_p_miso),
	.IOB(sampler6_adc_spi_n_miso),
	.O(main_spimaster0_interface_miso1)
);

OBUFTDS OBUFTDS_11(
	.I(main_spimaster1_interface_cs3),
	.T(main_spimaster1_interface_offline1),
	.O(sampler6_pgia_spi_p_cs_n),
	.OB(sampler6_pgia_spi_n_cs_n)
);

OBUFTDS OBUFTDS_12(
	.I(main_spimaster1_interface_clk1),
	.T(main_spimaster1_interface_offline1),
	.O(sampler6_pgia_spi_p_clk),
	.OB(sampler6_pgia_spi_n_clk)
);

IOBUFDS IOBUFDS_27(
	.I(main_spimaster1_interface_sdo1),
	.T((main_spimaster1_interface_offline1 | main_spimaster1_interface_half_duplex1)),
	.IO(sampler6_pgia_spi_p_mosi),
	.IOB(sampler6_pgia_spi_n_mosi),
	.O(main_spimaster1_interface_mosi1)
);

IOBUFDS IOBUFDS_28(
	.I(main_spimaster1_interface_sdo1),
	.T(1'd1),
	.IO(sampler6_pgia_spi_p_miso),
	.IOB(sampler6_pgia_spi_n_miso),
	.O(main_spimaster1_interface_miso1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_71 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x20_o[0] ^ 1'd0)),
	.D2((main_output_8x20_o[1] ^ 1'd0)),
	.D3((main_output_8x20_o[2] ^ 1'd0)),
	.D4((main_output_8x20_o[3] ^ 1'd0)),
	.D5((main_output_8x20_o[4] ^ 1'd0)),
	.D6((main_output_8x20_o[5] ^ 1'd0)),
	.D7((main_output_8x20_o[6] ^ 1'd0)),
	.D8((main_output_8x20_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x20_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x20_ser_out),
	.TQ(main_output_8x20_t_out)
);

IOBUFDS IOBUFDS_29(
	.I(main_output_8x20_ser_out),
	.T(main_output_8x20_t_out),
	.IO(sampler6_cnv_p),
	.IOB(sampler6_cnv_n)
);

OBUFTDS OBUFTDS_13(
	.I(main_spimaster2_interface_cs1[0]),
	.T(main_spimaster2_interface_offline),
	.O(zotino8_spi_p_cs_n[0]),
	.OB(zotino8_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_14(
	.I(main_spimaster2_interface_cs1[1]),
	.T(main_spimaster2_interface_offline),
	.O(zotino8_spi_p_cs_n[1]),
	.OB(zotino8_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_15(
	.I(main_spimaster2_interface_clk),
	.T(main_spimaster2_interface_offline),
	.O(zotino8_spi_p_clk),
	.OB(zotino8_spi_n_clk)
);

IOBUFDS IOBUFDS_30(
	.I(main_spimaster2_interface_sdo),
	.T((main_spimaster2_interface_offline | main_spimaster2_interface_half_duplex)),
	.IO(zotino8_spi_p_mosi),
	.IOB(zotino8_spi_n_mosi),
	.O(main_spimaster2_interface_mosi)
);

IOBUFDS IOBUFDS_31(
	.I(main_spimaster2_interface_sdo),
	.T(1'd1),
	.IO(zotino8_spi_p_miso),
	.IOB(zotino8_spi_n_miso),
	.O(main_spimaster2_interface_miso)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_72 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_ldac_phy_o[0] ^ 1'd0)),
	.D2((main_ldac_phy_o[1] ^ 1'd0)),
	.D3((main_ldac_phy_o[2] ^ 1'd0)),
	.D4((main_ldac_phy_o[3] ^ 1'd0)),
	.D5((main_ldac_phy_o[4] ^ 1'd0)),
	.D6((main_ldac_phy_o[5] ^ 1'd0)),
	.D7((main_ldac_phy_o[6] ^ 1'd0)),
	.D8((main_ldac_phy_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_ldac_phy_t_in),
	.TCE(1'd1),
	.OQ(main_ldac_phy_ser_out),
	.TQ(main_ldac_phy_t_out)
);

IOBUFDS IOBUFDS_32(
	.I(main_ldac_phy_ser_out),
	.T(main_ldac_phy_t_out),
	.IO(zotino8_ldac_n_p),
	.IOB(zotino8_ldac_n_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_73 (
	.CLK(sys4x_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_clr_phy_o[0] ^ 1'd0)),
	.D2((main_clr_phy_o[1] ^ 1'd0)),
	.D3((main_clr_phy_o[2] ^ 1'd0)),
	.D4((main_clr_phy_o[3] ^ 1'd0)),
	.D5((main_clr_phy_o[4] ^ 1'd0)),
	.D6((main_clr_phy_o[5] ^ 1'd0)),
	.D7((main_clr_phy_o[6] ^ 1'd0)),
	.D8((main_clr_phy_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_clr_phy_t_in),
	.TCE(1'd1),
	.OQ(main_clr_phy_ser_out),
	.TQ(main_clr_phy_t_out)
);

IOBUFDS IOBUFDS_33(
	.I(main_clr_phy_ser_out),
	.T(main_clr_phy_t_out),
	.IO(zotino8_clr_n_p),
	.IOB(zotino8_clr_n_n)
);

reg [13:0] latency_compensation[0:37];
reg [5:0] memadr_15;
always @(posedge rio_clk) begin : mem_write_block_25
	memadr_15 <= main_genericstandalone_rtio_core_sed_lane_dist_adr;
end

assign main_genericstandalone_rtio_core_sed_lane_dist_dat_r = latency_compensation[memadr_15];

initial begin
	$readmemh("latency_compensation.init", latency_compensation);
end

reg [116:0] storage_7[0:127];
reg [116:0] memdat_5;
reg [116:0] memdat_6;
always @(posedge rio_clk) begin : mem_write_block_26
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_we)
		storage_7[main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_dat_w;
	memdat_5 <= storage_7[main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_27
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_re)
		memdat_6 <= storage_7[main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_wrport_dat_r = memdat_5;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered0_rdport_dat_r = memdat_6;

reg [116:0] storage_8[0:127];
reg [116:0] memdat_7;
reg [116:0] memdat_8;
always @(posedge rio_clk) begin : mem_write_block_28
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_we)
		storage_8[main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_dat_w;
	memdat_7 <= storage_8[main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_29
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_re)
		memdat_8 <= storage_8[main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_wrport_dat_r = memdat_7;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered1_rdport_dat_r = memdat_8;

reg [116:0] storage_9[0:127];
reg [116:0] memdat_9;
reg [116:0] memdat_10;
always @(posedge rio_clk) begin : mem_write_block_30
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_we)
		storage_9[main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_dat_w;
	memdat_9 <= storage_9[main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_31
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_re)
		memdat_10 <= storage_9[main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_wrport_dat_r = memdat_9;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered2_rdport_dat_r = memdat_10;

reg [116:0] storage_10[0:127];
reg [116:0] memdat_11;
reg [116:0] memdat_12;
always @(posedge rio_clk) begin : mem_write_block_32
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_we)
		storage_10[main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_dat_w;
	memdat_11 <= storage_10[main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_33
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_re)
		memdat_12 <= storage_10[main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_wrport_dat_r = memdat_11;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered3_rdport_dat_r = memdat_12;

reg [116:0] storage_11[0:127];
reg [116:0] memdat_13;
reg [116:0] memdat_14;
always @(posedge rio_clk) begin : mem_write_block_34
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_we)
		storage_11[main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_dat_w;
	memdat_13 <= storage_11[main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_35
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_re)
		memdat_14 <= storage_11[main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_wrport_dat_r = memdat_13;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered4_rdport_dat_r = memdat_14;

reg [116:0] storage_12[0:127];
reg [116:0] memdat_15;
reg [116:0] memdat_16;
always @(posedge rio_clk) begin : mem_write_block_36
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_we)
		storage_12[main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_dat_w;
	memdat_15 <= storage_12[main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_37
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_re)
		memdat_16 <= storage_12[main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_wrport_dat_r = memdat_15;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered5_rdport_dat_r = memdat_16;

reg [116:0] storage_13[0:127];
reg [116:0] memdat_17;
reg [116:0] memdat_18;
always @(posedge rio_clk) begin : mem_write_block_38
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_we)
		storage_13[main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_dat_w;
	memdat_17 <= storage_13[main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_39
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_re)
		memdat_18 <= storage_13[main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_wrport_dat_r = memdat_17;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered6_rdport_dat_r = memdat_18;

reg [116:0] storage_14[0:127];
reg [116:0] memdat_19;
reg [116:0] memdat_20;
always @(posedge rio_clk) begin : mem_write_block_40
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_we)
		storage_14[main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_dat_w;
	memdat_19 <= storage_14[main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_41
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_re)
		memdat_20 <= storage_14[main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_wrport_dat_r = memdat_19;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered7_rdport_dat_r = memdat_20;

reg [116:0] storage_15[0:127];
reg [116:0] memdat_21;
reg [116:0] memdat_22;
always @(posedge rio_clk) begin : mem_write_block_42
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_we)
		storage_15[main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_dat_w;
	memdat_21 <= storage_15[main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_43
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_re)
		memdat_22 <= storage_15[main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_wrport_dat_r = memdat_21;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered8_rdport_dat_r = memdat_22;

reg [116:0] storage_16[0:127];
reg [116:0] memdat_23;
reg [116:0] memdat_24;
always @(posedge rio_clk) begin : mem_write_block_44
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_we)
		storage_16[main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_dat_w;
	memdat_23 <= storage_16[main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_45
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_re)
		memdat_24 <= storage_16[main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_wrport_dat_r = memdat_23;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered9_rdport_dat_r = memdat_24;

reg [116:0] storage_17[0:127];
reg [116:0] memdat_25;
reg [116:0] memdat_26;
always @(posedge rio_clk) begin : mem_write_block_46
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_we)
		storage_17[main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_dat_w;
	memdat_25 <= storage_17[main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_47
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_re)
		memdat_26 <= storage_17[main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_wrport_dat_r = memdat_25;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered10_rdport_dat_r = memdat_26;

reg [116:0] storage_18[0:127];
reg [116:0] memdat_27;
reg [116:0] memdat_28;
always @(posedge rio_clk) begin : mem_write_block_48
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_we)
		storage_18[main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_dat_w;
	memdat_27 <= storage_18[main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_49
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_re)
		memdat_28 <= storage_18[main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_wrport_dat_r = memdat_27;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered11_rdport_dat_r = memdat_28;

reg [116:0] storage_19[0:127];
reg [116:0] memdat_29;
reg [116:0] memdat_30;
always @(posedge rio_clk) begin : mem_write_block_50
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_we)
		storage_19[main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_dat_w;
	memdat_29 <= storage_19[main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_51
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_re)
		memdat_30 <= storage_19[main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_wrport_dat_r = memdat_29;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered12_rdport_dat_r = memdat_30;

reg [116:0] storage_20[0:127];
reg [116:0] memdat_31;
reg [116:0] memdat_32;
always @(posedge rio_clk) begin : mem_write_block_52
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_we)
		storage_20[main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_dat_w;
	memdat_31 <= storage_20[main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_53
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_re)
		memdat_32 <= storage_20[main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_wrport_dat_r = memdat_31;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered13_rdport_dat_r = memdat_32;

reg [116:0] storage_21[0:127];
reg [116:0] memdat_33;
reg [116:0] memdat_34;
always @(posedge rio_clk) begin : mem_write_block_54
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_we)
		storage_21[main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_dat_w;
	memdat_33 <= storage_21[main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_55
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_re)
		memdat_34 <= storage_21[main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_wrport_dat_r = memdat_33;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered14_rdport_dat_r = memdat_34;

reg [116:0] storage_22[0:127];
reg [116:0] memdat_35;
reg [116:0] memdat_36;
always @(posedge rio_clk) begin : mem_write_block_56
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_we)
		storage_22[main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_adr] <= main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_dat_w;
	memdat_35 <= storage_22[main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_57
	if (main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_re)
		memdat_36 <= storage_22[main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_adr];
end

assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_wrport_dat_r = memdat_35;
assign main_genericstandalone_rtio_core_sed_syncfifobuffered15_rdport_dat_r = memdat_36;

reg [0:0] en_replaces_rom[0:37];
reg [5:0] memadr_16;
always @(posedge rio_clk) begin : mem_write_block_58
	memadr_16 <= main_genericstandalone_rtio_core_sed_memory0_adr;
end

assign main_genericstandalone_rtio_core_sed_memory0_dat_r = en_replaces_rom[memadr_16];

initial begin
	$readmemh("en_replaces_rom.init", en_replaces_rom);
end

reg [0:0] en_replaces_rom_1[0:37];
reg [5:0] memadr_17;
always @(posedge rio_clk) begin : mem_write_block_59
	memadr_17 <= main_genericstandalone_rtio_core_sed_memory1_adr;
end

assign main_genericstandalone_rtio_core_sed_memory1_dat_r = en_replaces_rom_1[memadr_17];

initial begin
	$readmemh("en_replaces_rom_1.init", en_replaces_rom_1);
end

reg [0:0] en_replaces_rom_2[0:37];
reg [5:0] memadr_18;
always @(posedge rio_clk) begin : mem_write_block_60
	memadr_18 <= main_genericstandalone_rtio_core_sed_memory2_adr;
end

assign main_genericstandalone_rtio_core_sed_memory2_dat_r = en_replaces_rom_2[memadr_18];

initial begin
	$readmemh("en_replaces_rom_2.init", en_replaces_rom_2);
end

reg [0:0] en_replaces_rom_3[0:37];
reg [5:0] memadr_19;
always @(posedge rio_clk) begin : mem_write_block_61
	memadr_19 <= main_genericstandalone_rtio_core_sed_memory3_adr;
end

assign main_genericstandalone_rtio_core_sed_memory3_dat_r = en_replaces_rom_3[memadr_19];

initial begin
	$readmemh("en_replaces_rom_3.init", en_replaces_rom_3);
end

reg [0:0] en_replaces_rom_4[0:37];
reg [5:0] memadr_20;
always @(posedge rio_clk) begin : mem_write_block_62
	memadr_20 <= main_genericstandalone_rtio_core_sed_memory4_adr;
end

assign main_genericstandalone_rtio_core_sed_memory4_dat_r = en_replaces_rom_4[memadr_20];

initial begin
	$readmemh("en_replaces_rom_4.init", en_replaces_rom_4);
end

reg [0:0] en_replaces_rom_5[0:37];
reg [5:0] memadr_21;
always @(posedge rio_clk) begin : mem_write_block_63
	memadr_21 <= main_genericstandalone_rtio_core_sed_memory5_adr;
end

assign main_genericstandalone_rtio_core_sed_memory5_dat_r = en_replaces_rom_5[memadr_21];

initial begin
	$readmemh("en_replaces_rom_5.init", en_replaces_rom_5);
end

reg [0:0] en_replaces_rom_6[0:37];
reg [5:0] memadr_22;
always @(posedge rio_clk) begin : mem_write_block_64
	memadr_22 <= main_genericstandalone_rtio_core_sed_memory6_adr;
end

assign main_genericstandalone_rtio_core_sed_memory6_dat_r = en_replaces_rom_6[memadr_22];

initial begin
	$readmemh("en_replaces_rom_6.init", en_replaces_rom_6);
end

reg [0:0] en_replaces_rom_7[0:37];
reg [5:0] memadr_23;
always @(posedge rio_clk) begin : mem_write_block_65
	memadr_23 <= main_genericstandalone_rtio_core_sed_memory7_adr;
end

assign main_genericstandalone_rtio_core_sed_memory7_dat_r = en_replaces_rom_7[memadr_23];

initial begin
	$readmemh("en_replaces_rom_7.init", en_replaces_rom_7);
end

reg [0:0] en_replaces_rom_8[0:37];
reg [5:0] memadr_24;
always @(posedge rio_clk) begin : mem_write_block_66
	memadr_24 <= main_genericstandalone_rtio_core_sed_memory8_adr;
end

assign main_genericstandalone_rtio_core_sed_memory8_dat_r = en_replaces_rom_8[memadr_24];

initial begin
	$readmemh("en_replaces_rom_8.init", en_replaces_rom_8);
end

reg [0:0] en_replaces_rom_9[0:37];
reg [5:0] memadr_25;
always @(posedge rio_clk) begin : mem_write_block_67
	memadr_25 <= main_genericstandalone_rtio_core_sed_memory9_adr;
end

assign main_genericstandalone_rtio_core_sed_memory9_dat_r = en_replaces_rom_9[memadr_25];

initial begin
	$readmemh("en_replaces_rom_9.init", en_replaces_rom_9);
end

reg [0:0] en_replaces_rom_10[0:37];
reg [5:0] memadr_26;
always @(posedge rio_clk) begin : mem_write_block_68
	memadr_26 <= main_genericstandalone_rtio_core_sed_memory10_adr;
end

assign main_genericstandalone_rtio_core_sed_memory10_dat_r = en_replaces_rom_10[memadr_26];

initial begin
	$readmemh("en_replaces_rom_10.init", en_replaces_rom_10);
end

reg [0:0] en_replaces_rom_11[0:37];
reg [5:0] memadr_27;
always @(posedge rio_clk) begin : mem_write_block_69
	memadr_27 <= main_genericstandalone_rtio_core_sed_memory11_adr;
end

assign main_genericstandalone_rtio_core_sed_memory11_dat_r = en_replaces_rom_11[memadr_27];

initial begin
	$readmemh("en_replaces_rom_11.init", en_replaces_rom_11);
end

reg [0:0] en_replaces_rom_12[0:37];
reg [5:0] memadr_28;
always @(posedge rio_clk) begin : mem_write_block_70
	memadr_28 <= main_genericstandalone_rtio_core_sed_memory12_adr;
end

assign main_genericstandalone_rtio_core_sed_memory12_dat_r = en_replaces_rom_12[memadr_28];

initial begin
	$readmemh("en_replaces_rom_12.init", en_replaces_rom_12);
end

reg [0:0] en_replaces_rom_13[0:37];
reg [5:0] memadr_29;
always @(posedge rio_clk) begin : mem_write_block_71
	memadr_29 <= main_genericstandalone_rtio_core_sed_memory13_adr;
end

assign main_genericstandalone_rtio_core_sed_memory13_dat_r = en_replaces_rom_13[memadr_29];

initial begin
	$readmemh("en_replaces_rom_13.init", en_replaces_rom_13);
end

reg [0:0] en_replaces_rom_14[0:37];
reg [5:0] memadr_30;
always @(posedge rio_clk) begin : mem_write_block_72
	memadr_30 <= main_genericstandalone_rtio_core_sed_memory14_adr;
end

assign main_genericstandalone_rtio_core_sed_memory14_dat_r = en_replaces_rom_14[memadr_30];

initial begin
	$readmemh("en_replaces_rom_14.init", en_replaces_rom_14);
end

reg [0:0] en_replaces_rom_15[0:37];
reg [5:0] memadr_31;
always @(posedge rio_clk) begin : mem_write_block_73
	memadr_31 <= main_genericstandalone_rtio_core_sed_memory15_adr;
end

assign main_genericstandalone_rtio_core_sed_memory15_dat_r = en_replaces_rom_15[memadr_31];

initial begin
	$readmemh("en_replaces_rom_15.init", en_replaces_rom_15);
end

reg [64:0] storage_23[0:63];
reg [64:0] memdat_37;
reg [64:0] memdat_38;
always @(posedge rio_clk) begin : mem_write_block_74
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_we)
		storage_23[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_dat_w;
	memdat_37 <= storage_23[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_75
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_re)
		memdat_38 <= storage_23[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_wrport_dat_r = memdat_37;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered0_rdport_dat_r = memdat_38;

reg [64:0] storage_24[0:63];
reg [64:0] memdat_39;
reg [64:0] memdat_40;
always @(posedge rio_clk) begin : mem_write_block_76
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_we)
		storage_24[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_dat_w;
	memdat_39 <= storage_24[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_77
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_re)
		memdat_40 <= storage_24[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_wrport_dat_r = memdat_39;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered1_rdport_dat_r = memdat_40;

reg [64:0] storage_25[0:63];
reg [64:0] memdat_41;
reg [64:0] memdat_42;
always @(posedge rio_clk) begin : mem_write_block_78
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_we)
		storage_25[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_dat_w;
	memdat_41 <= storage_25[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_79
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_re)
		memdat_42 <= storage_25[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_wrport_dat_r = memdat_41;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered2_rdport_dat_r = memdat_42;

reg [64:0] storage_26[0:63];
reg [64:0] memdat_43;
reg [64:0] memdat_44;
always @(posedge rio_clk) begin : mem_write_block_80
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_we)
		storage_26[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_dat_w;
	memdat_43 <= storage_26[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_81
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_re)
		memdat_44 <= storage_26[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_wrport_dat_r = memdat_43;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered3_rdport_dat_r = memdat_44;

reg [31:0] storage_27[0:3];
reg [31:0] memdat_45;
reg [31:0] memdat_46;
always @(posedge rio_clk) begin : mem_write_block_82
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_we)
		storage_27[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_dat_w;
	memdat_45 <= storage_27[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_83
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_re)
		memdat_46 <= storage_27[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_wrport_dat_r = memdat_45;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered4_rdport_dat_r = memdat_46;

reg [31:0] storage_28[0:3];
reg [31:0] memdat_47;
reg [31:0] memdat_48;
always @(posedge rio_clk) begin : mem_write_block_84
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_we)
		storage_28[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_dat_w;
	memdat_47 <= storage_28[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_85
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_re)
		memdat_48 <= storage_28[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_wrport_dat_r = memdat_47;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered5_rdport_dat_r = memdat_48;

reg [31:0] storage_29[0:3];
reg [31:0] memdat_49;
reg [31:0] memdat_50;
always @(posedge rio_clk) begin : mem_write_block_86
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_we)
		storage_29[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_dat_w;
	memdat_49 <= storage_29[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_87
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_re)
		memdat_50 <= storage_29[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_wrport_dat_r = memdat_49;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered6_rdport_dat_r = memdat_50;

reg [31:0] storage_30[0:3];
reg [31:0] memdat_51;
reg [31:0] memdat_52;
always @(posedge rio_clk) begin : mem_write_block_88
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_we)
		storage_30[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_dat_w;
	memdat_51 <= storage_30[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_89
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_re)
		memdat_52 <= storage_30[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_wrport_dat_r = memdat_51;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered7_rdport_dat_r = memdat_52;

reg [31:0] storage_31[0:3];
reg [31:0] memdat_53;
reg [31:0] memdat_54;
always @(posedge rio_clk) begin : mem_write_block_90
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_we)
		storage_31[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_adr] <= main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_dat_w;
	memdat_53 <= storage_31[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_adr];
end

always @(posedge rio_clk) begin : mem_write_block_91
	if (main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_re)
		memdat_54 <= storage_31[main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_adr];
end

assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_wrport_dat_r = memdat_53;
assign main_genericstandalone_rtio_core_inputcollector_syncfifobuffered8_rdport_dat_r = memdat_54;

reg [128:0] storage_32[0:127];
reg [128:0] memdat_55;
reg [128:0] memdat_56;
always @(posedge sys_kernel_clk) begin : mem_write_block_92
	if (main_genericstandalone_dma_fifo_wrport_we)
		storage_32[main_genericstandalone_dma_fifo_wrport_adr] <= main_genericstandalone_dma_fifo_wrport_dat_w;
	memdat_55 <= storage_32[main_genericstandalone_dma_fifo_wrport_adr];
end

always @(posedge sys_kernel_clk) begin : mem_write_block_93
	if (main_genericstandalone_dma_fifo_rdport_re)
		memdat_56 <= storage_32[main_genericstandalone_dma_fifo_rdport_adr];
end

assign main_genericstandalone_dma_fifo_wrport_dat_r = memdat_55;
assign main_genericstandalone_dma_fifo_rdport_dat_r = memdat_56;

reg [256:0] storage_33[0:127];
reg [256:0] memdat_57;
reg [256:0] memdat_58;
always @(posedge sys_clk) begin : mem_write_block_94
	if (main_genericstandalone_rtio_analyzer_fifo_wrport_we)
		storage_33[main_genericstandalone_rtio_analyzer_fifo_wrport_adr] <= main_genericstandalone_rtio_analyzer_fifo_wrport_dat_w;
	memdat_57 <= storage_33[main_genericstandalone_rtio_analyzer_fifo_wrport_adr];
end

always @(posedge sys_clk) begin : mem_write_block_95
	if (main_genericstandalone_rtio_analyzer_fifo_rdport_re)
		memdat_58 <= storage_33[main_genericstandalone_rtio_analyzer_fifo_rdport_adr];
end

assign main_genericstandalone_rtio_analyzer_fifo_wrport_dat_r = memdat_57;
assign main_genericstandalone_rtio_analyzer_fifo_rdport_dat_r = memdat_58;

reg [7:0] mem_grain0[0:190];
reg [7:0] memadr_32;
reg [7:0] memadr_33;
always @(posedge sys_clk) begin : mem_write_block_96
	memadr_32 <= main_genericstandalone_sram158_adr;
end

always @(posedge sys_clk) begin : mem_write_block_97
	if (main_genericstandalone_sram4_we[0])
		mem_grain0[main_genericstandalone_sram4_adr] <= main_genericstandalone_sram4_dat_w[7:0];
	memadr_33 <= main_genericstandalone_sram4_adr;
end

assign main_genericstandalone_sram159_dat_r[7:0] = mem_grain0[memadr_32];
assign main_genericstandalone_sram4_dat_r[7:0] = mem_grain0[memadr_33];

reg [7:0] mem_grain1[0:190];
reg [7:0] memadr_34;
reg [7:0] memadr_35;
always @(posedge sys_clk) begin : mem_write_block_98
	memadr_34 <= main_genericstandalone_sram158_adr;
end

always @(posedge sys_clk) begin : mem_write_block_99
	if (main_genericstandalone_sram4_we[1])
		mem_grain1[main_genericstandalone_sram4_adr] <= main_genericstandalone_sram4_dat_w[15:8];
	memadr_35 <= main_genericstandalone_sram4_adr;
end

assign main_genericstandalone_sram159_dat_r[15:8] = mem_grain1[memadr_34];
assign main_genericstandalone_sram4_dat_r[15:8] = mem_grain1[memadr_35];

reg [7:0] mem_grain2[0:190];
reg [7:0] memadr_36;
reg [7:0] memadr_37;
always @(posedge sys_clk) begin : mem_write_block_100
	memadr_36 <= main_genericstandalone_sram158_adr;
end

always @(posedge sys_clk) begin : mem_write_block_101
	if (main_genericstandalone_sram4_we[2])
		mem_grain2[main_genericstandalone_sram4_adr] <= main_genericstandalone_sram4_dat_w[23:16];
	memadr_37 <= main_genericstandalone_sram4_adr;
end

assign main_genericstandalone_sram159_dat_r[23:16] = mem_grain2[memadr_36];
assign main_genericstandalone_sram4_dat_r[23:16] = mem_grain2[memadr_37];

reg [7:0] mem_grain3[0:190];
reg [7:0] memadr_38;
reg [7:0] memadr_39;
always @(posedge sys_clk) begin : mem_write_block_102
	memadr_38 <= main_genericstandalone_sram158_adr;
end

always @(posedge sys_clk) begin : mem_write_block_103
	if (main_genericstandalone_sram4_we[3])
		mem_grain3[main_genericstandalone_sram4_adr] <= main_genericstandalone_sram4_dat_w[31:24];
	memadr_39 <= main_genericstandalone_sram4_adr;
end

assign main_genericstandalone_sram159_dat_r[31:24] = mem_grain3[memadr_38];
assign main_genericstandalone_sram4_dat_r[31:24] = mem_grain3[memadr_39];

reg [7:0] mem_grain4[0:190];
reg [7:0] memadr_40;
reg [7:0] memadr_41;
always @(posedge sys_clk) begin : mem_write_block_104
	memadr_40 <= main_genericstandalone_sram158_adr;
end

always @(posedge sys_clk) begin : mem_write_block_105
	if (main_genericstandalone_sram4_we[4])
		mem_grain4[main_genericstandalone_sram4_adr] <= main_genericstandalone_sram4_dat_w[39:32];
	memadr_41 <= main_genericstandalone_sram4_adr;
end

assign main_genericstandalone_sram159_dat_r[39:32] = mem_grain4[memadr_40];
assign main_genericstandalone_sram4_dat_r[39:32] = mem_grain4[memadr_41];

reg [7:0] mem_grain5[0:190];
reg [7:0] memadr_42;
reg [7:0] memadr_43;
always @(posedge sys_clk) begin : mem_write_block_106
	memadr_42 <= main_genericstandalone_sram158_adr;
end

always @(posedge sys_clk) begin : mem_write_block_107
	if (main_genericstandalone_sram4_we[5])
		mem_grain5[main_genericstandalone_sram4_adr] <= main_genericstandalone_sram4_dat_w[47:40];
	memadr_43 <= main_genericstandalone_sram4_adr;
end

assign main_genericstandalone_sram159_dat_r[47:40] = mem_grain5[memadr_42];
assign main_genericstandalone_sram4_dat_r[47:40] = mem_grain5[memadr_43];

reg [7:0] mem_grain6[0:190];
reg [7:0] memadr_44;
reg [7:0] memadr_45;
always @(posedge sys_clk) begin : mem_write_block_108
	memadr_44 <= main_genericstandalone_sram158_adr;
end

always @(posedge sys_clk) begin : mem_write_block_109
	if (main_genericstandalone_sram4_we[6])
		mem_grain6[main_genericstandalone_sram4_adr] <= main_genericstandalone_sram4_dat_w[55:48];
	memadr_45 <= main_genericstandalone_sram4_adr;
end

assign main_genericstandalone_sram159_dat_r[55:48] = mem_grain6[memadr_44];
assign main_genericstandalone_sram4_dat_r[55:48] = mem_grain6[memadr_45];

reg [7:0] mem_grain7[0:190];
reg [7:0] memadr_46;
reg [7:0] memadr_47;
always @(posedge sys_clk) begin : mem_write_block_110
	memadr_46 <= main_genericstandalone_sram158_adr;
end

always @(posedge sys_clk) begin : mem_write_block_111
	if (main_genericstandalone_sram4_we[7])
		mem_grain7[main_genericstandalone_sram4_adr] <= main_genericstandalone_sram4_dat_w[63:56];
	memadr_47 <= main_genericstandalone_sram4_adr;
end

assign main_genericstandalone_sram159_dat_r[63:56] = mem_grain7[memadr_46];
assign main_genericstandalone_sram4_dat_r[63:56] = mem_grain7[memadr_47];

reg [7:0] mem_grain0_1[0:190];
reg [7:0] memadr_48;
reg [7:0] memadr_49;
always @(posedge sys_clk) begin : mem_write_block_112
	memadr_48 <= main_genericstandalone_sram160_adr;
end

always @(posedge sys_clk) begin : mem_write_block_113
	if (main_genericstandalone_sram5_we[0])
		mem_grain0_1[main_genericstandalone_sram5_adr] <= main_genericstandalone_sram5_dat_w[7:0];
	memadr_49 <= main_genericstandalone_sram5_adr;
end

assign main_genericstandalone_sram161_dat_r[7:0] = mem_grain0_1[memadr_48];
assign main_genericstandalone_sram5_dat_r[7:0] = mem_grain0_1[memadr_49];

reg [7:0] mem_grain1_1[0:190];
reg [7:0] memadr_50;
reg [7:0] memadr_51;
always @(posedge sys_clk) begin : mem_write_block_114
	memadr_50 <= main_genericstandalone_sram160_adr;
end

always @(posedge sys_clk) begin : mem_write_block_115
	if (main_genericstandalone_sram5_we[1])
		mem_grain1_1[main_genericstandalone_sram5_adr] <= main_genericstandalone_sram5_dat_w[15:8];
	memadr_51 <= main_genericstandalone_sram5_adr;
end

assign main_genericstandalone_sram161_dat_r[15:8] = mem_grain1_1[memadr_50];
assign main_genericstandalone_sram5_dat_r[15:8] = mem_grain1_1[memadr_51];

reg [7:0] mem_grain2_1[0:190];
reg [7:0] memadr_52;
reg [7:0] memadr_53;
always @(posedge sys_clk) begin : mem_write_block_116
	memadr_52 <= main_genericstandalone_sram160_adr;
end

always @(posedge sys_clk) begin : mem_write_block_117
	if (main_genericstandalone_sram5_we[2])
		mem_grain2_1[main_genericstandalone_sram5_adr] <= main_genericstandalone_sram5_dat_w[23:16];
	memadr_53 <= main_genericstandalone_sram5_adr;
end

assign main_genericstandalone_sram161_dat_r[23:16] = mem_grain2_1[memadr_52];
assign main_genericstandalone_sram5_dat_r[23:16] = mem_grain2_1[memadr_53];

reg [7:0] mem_grain3_1[0:190];
reg [7:0] memadr_54;
reg [7:0] memadr_55;
always @(posedge sys_clk) begin : mem_write_block_118
	memadr_54 <= main_genericstandalone_sram160_adr;
end

always @(posedge sys_clk) begin : mem_write_block_119
	if (main_genericstandalone_sram5_we[3])
		mem_grain3_1[main_genericstandalone_sram5_adr] <= main_genericstandalone_sram5_dat_w[31:24];
	memadr_55 <= main_genericstandalone_sram5_adr;
end

assign main_genericstandalone_sram161_dat_r[31:24] = mem_grain3_1[memadr_54];
assign main_genericstandalone_sram5_dat_r[31:24] = mem_grain3_1[memadr_55];

reg [7:0] mem_grain4_1[0:190];
reg [7:0] memadr_56;
reg [7:0] memadr_57;
always @(posedge sys_clk) begin : mem_write_block_120
	memadr_56 <= main_genericstandalone_sram160_adr;
end

always @(posedge sys_clk) begin : mem_write_block_121
	if (main_genericstandalone_sram5_we[4])
		mem_grain4_1[main_genericstandalone_sram5_adr] <= main_genericstandalone_sram5_dat_w[39:32];
	memadr_57 <= main_genericstandalone_sram5_adr;
end

assign main_genericstandalone_sram161_dat_r[39:32] = mem_grain4_1[memadr_56];
assign main_genericstandalone_sram5_dat_r[39:32] = mem_grain4_1[memadr_57];

reg [7:0] mem_grain5_1[0:190];
reg [7:0] memadr_58;
reg [7:0] memadr_59;
always @(posedge sys_clk) begin : mem_write_block_122
	memadr_58 <= main_genericstandalone_sram160_adr;
end

always @(posedge sys_clk) begin : mem_write_block_123
	if (main_genericstandalone_sram5_we[5])
		mem_grain5_1[main_genericstandalone_sram5_adr] <= main_genericstandalone_sram5_dat_w[47:40];
	memadr_59 <= main_genericstandalone_sram5_adr;
end

assign main_genericstandalone_sram161_dat_r[47:40] = mem_grain5_1[memadr_58];
assign main_genericstandalone_sram5_dat_r[47:40] = mem_grain5_1[memadr_59];

reg [7:0] mem_grain6_1[0:190];
reg [7:0] memadr_60;
reg [7:0] memadr_61;
always @(posedge sys_clk) begin : mem_write_block_124
	memadr_60 <= main_genericstandalone_sram160_adr;
end

always @(posedge sys_clk) begin : mem_write_block_125
	if (main_genericstandalone_sram5_we[6])
		mem_grain6_1[main_genericstandalone_sram5_adr] <= main_genericstandalone_sram5_dat_w[55:48];
	memadr_61 <= main_genericstandalone_sram5_adr;
end

assign main_genericstandalone_sram161_dat_r[55:48] = mem_grain6_1[memadr_60];
assign main_genericstandalone_sram5_dat_r[55:48] = mem_grain6_1[memadr_61];

reg [7:0] mem_grain7_1[0:190];
reg [7:0] memadr_62;
reg [7:0] memadr_63;
always @(posedge sys_clk) begin : mem_write_block_126
	memadr_62 <= main_genericstandalone_sram160_adr;
end

always @(posedge sys_clk) begin : mem_write_block_127
	if (main_genericstandalone_sram5_we[7])
		mem_grain7_1[main_genericstandalone_sram5_adr] <= main_genericstandalone_sram5_dat_w[63:56];
	memadr_63 <= main_genericstandalone_sram5_adr;
end

assign main_genericstandalone_sram161_dat_r[63:56] = mem_grain7_1[memadr_62];
assign main_genericstandalone_sram5_dat_r[63:56] = mem_grain7_1[memadr_63];

reg [7:0] mem_grain0_2[0:190];
reg [7:0] memadr_64;
reg [7:0] memadr_65;
always @(posedge sys_clk) begin : mem_write_block_128
	memadr_64 <= main_genericstandalone_sram162_adr;
end

always @(posedge sys_clk) begin : mem_write_block_129
	if (main_genericstandalone_sram6_we[0])
		mem_grain0_2[main_genericstandalone_sram6_adr] <= main_genericstandalone_sram6_dat_w[7:0];
	memadr_65 <= main_genericstandalone_sram6_adr;
end

assign main_genericstandalone_sram163_dat_r[7:0] = mem_grain0_2[memadr_64];
assign main_genericstandalone_sram6_dat_r[7:0] = mem_grain0_2[memadr_65];

reg [7:0] mem_grain1_2[0:190];
reg [7:0] memadr_66;
reg [7:0] memadr_67;
always @(posedge sys_clk) begin : mem_write_block_130
	memadr_66 <= main_genericstandalone_sram162_adr;
end

always @(posedge sys_clk) begin : mem_write_block_131
	if (main_genericstandalone_sram6_we[1])
		mem_grain1_2[main_genericstandalone_sram6_adr] <= main_genericstandalone_sram6_dat_w[15:8];
	memadr_67 <= main_genericstandalone_sram6_adr;
end

assign main_genericstandalone_sram163_dat_r[15:8] = mem_grain1_2[memadr_66];
assign main_genericstandalone_sram6_dat_r[15:8] = mem_grain1_2[memadr_67];

reg [7:0] mem_grain2_2[0:190];
reg [7:0] memadr_68;
reg [7:0] memadr_69;
always @(posedge sys_clk) begin : mem_write_block_132
	memadr_68 <= main_genericstandalone_sram162_adr;
end

always @(posedge sys_clk) begin : mem_write_block_133
	if (main_genericstandalone_sram6_we[2])
		mem_grain2_2[main_genericstandalone_sram6_adr] <= main_genericstandalone_sram6_dat_w[23:16];
	memadr_69 <= main_genericstandalone_sram6_adr;
end

assign main_genericstandalone_sram163_dat_r[23:16] = mem_grain2_2[memadr_68];
assign main_genericstandalone_sram6_dat_r[23:16] = mem_grain2_2[memadr_69];

reg [7:0] mem_grain3_2[0:190];
reg [7:0] memadr_70;
reg [7:0] memadr_71;
always @(posedge sys_clk) begin : mem_write_block_134
	memadr_70 <= main_genericstandalone_sram162_adr;
end

always @(posedge sys_clk) begin : mem_write_block_135
	if (main_genericstandalone_sram6_we[3])
		mem_grain3_2[main_genericstandalone_sram6_adr] <= main_genericstandalone_sram6_dat_w[31:24];
	memadr_71 <= main_genericstandalone_sram6_adr;
end

assign main_genericstandalone_sram163_dat_r[31:24] = mem_grain3_2[memadr_70];
assign main_genericstandalone_sram6_dat_r[31:24] = mem_grain3_2[memadr_71];

reg [7:0] mem_grain4_2[0:190];
reg [7:0] memadr_72;
reg [7:0] memadr_73;
always @(posedge sys_clk) begin : mem_write_block_136
	memadr_72 <= main_genericstandalone_sram162_adr;
end

always @(posedge sys_clk) begin : mem_write_block_137
	if (main_genericstandalone_sram6_we[4])
		mem_grain4_2[main_genericstandalone_sram6_adr] <= main_genericstandalone_sram6_dat_w[39:32];
	memadr_73 <= main_genericstandalone_sram6_adr;
end

assign main_genericstandalone_sram163_dat_r[39:32] = mem_grain4_2[memadr_72];
assign main_genericstandalone_sram6_dat_r[39:32] = mem_grain4_2[memadr_73];

reg [7:0] mem_grain5_2[0:190];
reg [7:0] memadr_74;
reg [7:0] memadr_75;
always @(posedge sys_clk) begin : mem_write_block_138
	memadr_74 <= main_genericstandalone_sram162_adr;
end

always @(posedge sys_clk) begin : mem_write_block_139
	if (main_genericstandalone_sram6_we[5])
		mem_grain5_2[main_genericstandalone_sram6_adr] <= main_genericstandalone_sram6_dat_w[47:40];
	memadr_75 <= main_genericstandalone_sram6_adr;
end

assign main_genericstandalone_sram163_dat_r[47:40] = mem_grain5_2[memadr_74];
assign main_genericstandalone_sram6_dat_r[47:40] = mem_grain5_2[memadr_75];

reg [7:0] mem_grain6_2[0:190];
reg [7:0] memadr_76;
reg [7:0] memadr_77;
always @(posedge sys_clk) begin : mem_write_block_140
	memadr_76 <= main_genericstandalone_sram162_adr;
end

always @(posedge sys_clk) begin : mem_write_block_141
	if (main_genericstandalone_sram6_we[6])
		mem_grain6_2[main_genericstandalone_sram6_adr] <= main_genericstandalone_sram6_dat_w[55:48];
	memadr_77 <= main_genericstandalone_sram6_adr;
end

assign main_genericstandalone_sram163_dat_r[55:48] = mem_grain6_2[memadr_76];
assign main_genericstandalone_sram6_dat_r[55:48] = mem_grain6_2[memadr_77];

reg [7:0] mem_grain7_2[0:190];
reg [7:0] memadr_78;
reg [7:0] memadr_79;
always @(posedge sys_clk) begin : mem_write_block_142
	memadr_78 <= main_genericstandalone_sram162_adr;
end

always @(posedge sys_clk) begin : mem_write_block_143
	if (main_genericstandalone_sram6_we[7])
		mem_grain7_2[main_genericstandalone_sram6_adr] <= main_genericstandalone_sram6_dat_w[63:56];
	memadr_79 <= main_genericstandalone_sram6_adr;
end

assign main_genericstandalone_sram163_dat_r[63:56] = mem_grain7_2[memadr_78];
assign main_genericstandalone_sram6_dat_r[63:56] = mem_grain7_2[memadr_79];

reg [7:0] mem_grain0_3[0:190];
reg [7:0] memadr_80;
reg [7:0] memadr_81;
always @(posedge sys_clk) begin : mem_write_block_144
	memadr_80 <= main_genericstandalone_sram164_adr;
end

always @(posedge sys_clk) begin : mem_write_block_145
	if (main_genericstandalone_sram7_we[0])
		mem_grain0_3[main_genericstandalone_sram7_adr] <= main_genericstandalone_sram7_dat_w[7:0];
	memadr_81 <= main_genericstandalone_sram7_adr;
end

assign main_genericstandalone_sram165_dat_r[7:0] = mem_grain0_3[memadr_80];
assign main_genericstandalone_sram7_dat_r[7:0] = mem_grain0_3[memadr_81];

reg [7:0] mem_grain1_3[0:190];
reg [7:0] memadr_82;
reg [7:0] memadr_83;
always @(posedge sys_clk) begin : mem_write_block_146
	memadr_82 <= main_genericstandalone_sram164_adr;
end

always @(posedge sys_clk) begin : mem_write_block_147
	if (main_genericstandalone_sram7_we[1])
		mem_grain1_3[main_genericstandalone_sram7_adr] <= main_genericstandalone_sram7_dat_w[15:8];
	memadr_83 <= main_genericstandalone_sram7_adr;
end

assign main_genericstandalone_sram165_dat_r[15:8] = mem_grain1_3[memadr_82];
assign main_genericstandalone_sram7_dat_r[15:8] = mem_grain1_3[memadr_83];

reg [7:0] mem_grain2_3[0:190];
reg [7:0] memadr_84;
reg [7:0] memadr_85;
always @(posedge sys_clk) begin : mem_write_block_148
	memadr_84 <= main_genericstandalone_sram164_adr;
end

always @(posedge sys_clk) begin : mem_write_block_149
	if (main_genericstandalone_sram7_we[2])
		mem_grain2_3[main_genericstandalone_sram7_adr] <= main_genericstandalone_sram7_dat_w[23:16];
	memadr_85 <= main_genericstandalone_sram7_adr;
end

assign main_genericstandalone_sram165_dat_r[23:16] = mem_grain2_3[memadr_84];
assign main_genericstandalone_sram7_dat_r[23:16] = mem_grain2_3[memadr_85];

reg [7:0] mem_grain3_3[0:190];
reg [7:0] memadr_86;
reg [7:0] memadr_87;
always @(posedge sys_clk) begin : mem_write_block_150
	memadr_86 <= main_genericstandalone_sram164_adr;
end

always @(posedge sys_clk) begin : mem_write_block_151
	if (main_genericstandalone_sram7_we[3])
		mem_grain3_3[main_genericstandalone_sram7_adr] <= main_genericstandalone_sram7_dat_w[31:24];
	memadr_87 <= main_genericstandalone_sram7_adr;
end

assign main_genericstandalone_sram165_dat_r[31:24] = mem_grain3_3[memadr_86];
assign main_genericstandalone_sram7_dat_r[31:24] = mem_grain3_3[memadr_87];

reg [7:0] mem_grain4_3[0:190];
reg [7:0] memadr_88;
reg [7:0] memadr_89;
always @(posedge sys_clk) begin : mem_write_block_152
	memadr_88 <= main_genericstandalone_sram164_adr;
end

always @(posedge sys_clk) begin : mem_write_block_153
	if (main_genericstandalone_sram7_we[4])
		mem_grain4_3[main_genericstandalone_sram7_adr] <= main_genericstandalone_sram7_dat_w[39:32];
	memadr_89 <= main_genericstandalone_sram7_adr;
end

assign main_genericstandalone_sram165_dat_r[39:32] = mem_grain4_3[memadr_88];
assign main_genericstandalone_sram7_dat_r[39:32] = mem_grain4_3[memadr_89];

reg [7:0] mem_grain5_3[0:190];
reg [7:0] memadr_90;
reg [7:0] memadr_91;
always @(posedge sys_clk) begin : mem_write_block_154
	memadr_90 <= main_genericstandalone_sram164_adr;
end

always @(posedge sys_clk) begin : mem_write_block_155
	if (main_genericstandalone_sram7_we[5])
		mem_grain5_3[main_genericstandalone_sram7_adr] <= main_genericstandalone_sram7_dat_w[47:40];
	memadr_91 <= main_genericstandalone_sram7_adr;
end

assign main_genericstandalone_sram165_dat_r[47:40] = mem_grain5_3[memadr_90];
assign main_genericstandalone_sram7_dat_r[47:40] = mem_grain5_3[memadr_91];

reg [7:0] mem_grain6_3[0:190];
reg [7:0] memadr_92;
reg [7:0] memadr_93;
always @(posedge sys_clk) begin : mem_write_block_156
	memadr_92 <= main_genericstandalone_sram164_adr;
end

always @(posedge sys_clk) begin : mem_write_block_157
	if (main_genericstandalone_sram7_we[6])
		mem_grain6_3[main_genericstandalone_sram7_adr] <= main_genericstandalone_sram7_dat_w[55:48];
	memadr_93 <= main_genericstandalone_sram7_adr;
end

assign main_genericstandalone_sram165_dat_r[55:48] = mem_grain6_3[memadr_92];
assign main_genericstandalone_sram7_dat_r[55:48] = mem_grain6_3[memadr_93];

reg [7:0] mem_grain7_3[0:190];
reg [7:0] memadr_94;
reg [7:0] memadr_95;
always @(posedge sys_clk) begin : mem_write_block_158
	memadr_94 <= main_genericstandalone_sram164_adr;
end

always @(posedge sys_clk) begin : mem_write_block_159
	if (main_genericstandalone_sram7_we[7])
		mem_grain7_3[main_genericstandalone_sram7_adr] <= main_genericstandalone_sram7_dat_w[63:56];
	memadr_95 <= main_genericstandalone_sram7_adr;
end

assign main_genericstandalone_sram165_dat_r[63:56] = mem_grain7_3[memadr_94];
assign main_genericstandalone_sram7_dat_r[63:56] = mem_grain7_3[memadr_95];

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl0_async_reset),
	.Q(builder_xilinxasyncresetsynchronizerimpl0_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl0_async_reset),
	.Q(clk200_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl1_async_reset),
	.Q(builder_xilinxasyncresetsynchronizerimpl1_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl1_async_reset),
	.Q(eth_tx_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl2_async_reset),
	.Q(builder_xilinxasyncresetsynchronizerimpl2_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl2_async_reset),
	.Q(eth_rx_rst)
);

OBUFDS OBUFDS_2(
	.I(1'd0),
	.O(urukul4_dds_reset_sync_in_p),
	.OB(urukul4_dds_reset_sync_in_n)
);

OBUFDS OBUFDS_3(
	.I(1'd1),
	.O(sampler6_sdr_p),
	.OB(sampler6_sdr_n)
);

endmodule
